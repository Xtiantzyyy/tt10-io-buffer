magic
tech sky130A
magscale 1 2
timestamp 1746118077
<< nwell >>
rect 21680 42270 23700 43400
rect 2399 42060 3039 42230
rect 21680 42150 23200 42270
rect 21680 42140 22150 42150
rect 2399 41450 3009 42060
rect 2399 40960 3089 41450
rect 3350 41020 5629 42040
rect 5909 41300 10019 42020
rect 3219 40230 4240 40720
rect 3219 39740 4239 40230
rect 4499 39740 5519 40720
rect 6309 39980 10009 40700
rect 15120 36260 24950 36410
rect 15120 35980 25400 36260
rect 15120 35680 16230 35980
rect 17300 35970 25400 35980
rect 17300 35770 21350 35970
rect 15120 35560 15680 35680
rect 17300 35530 20220 35770
rect 19260 34970 19510 35530
rect 20900 35520 21350 35770
rect 22300 35530 25400 35970
rect 20990 34980 21240 35520
rect 21000 34970 21240 34980
rect 24220 34970 24470 35530
rect 5390 34730 10920 34800
rect 3730 33930 10920 34730
rect 3730 33470 6330 33930
rect 13690 32310 14340 32570
rect 13690 32300 14338 32310
rect 13688 31830 14338 32300
rect 15990 31960 25450 32240
rect 17300 31870 25450 31960
rect 17300 31460 21410 31870
rect 22310 31460 25450 31870
rect 19260 30910 19780 31460
rect 21050 30920 21300 31460
rect 21060 30910 21300 30920
rect 24280 30900 24820 31460
rect 6310 30550 11300 30650
rect 3790 30480 11300 30550
rect 2130 29760 11300 30480
rect 2130 29220 6380 29760
rect 7270 25940 20680 26660
rect 7240 21610 20530 21630
rect 7240 20910 20680 21610
rect 7240 20070 8530 20520
rect 7240 19320 20680 20070
rect 9630 14250 21160 14950
rect 7240 12720 21160 13430
rect 7260 12710 8620 12720
rect 7800 10340 8430 10760
rect 7240 10330 9790 10340
rect 7240 9530 21160 10330
rect 9830 6880 17120 8300
rect 9810 4370 13280 5990
rect 13550 4620 17060 6040
<< pwell >>
rect 3640 37374 11100 37390
rect 3482 37088 11100 37374
rect 3640 35960 11100 37088
rect 7140 22720 20630 24860
rect 7050 17450 20730 18250
rect 19500 16780 20430 17450
<< nmos >>
rect 21790 41680 21820 41880
rect 23450 41900 23480 42100
rect 22650 41510 22680 41710
rect 22950 41510 22980 41710
rect 23060 41510 23090 41710
rect 23450 41370 23480 41570
rect 6019 40980 6049 41180
rect 6249 40980 6279 41180
rect 6359 40980 6389 41180
rect 6589 40980 6619 41180
rect 6699 40980 6729 41180
rect 6809 40980 6839 41180
rect 6919 40980 6949 41180
rect 7149 40980 7179 41180
rect 7259 40980 7289 41180
rect 7369 40980 7399 41180
rect 7479 40980 7509 41180
rect 7589 40980 7619 41180
rect 7699 40980 7729 41180
rect 7809 40980 7839 41180
rect 7919 40980 7949 41180
rect 8209 40980 8239 41180
rect 8319 40980 8349 41180
rect 8429 40980 8459 41180
rect 8539 40980 8569 41180
rect 8649 40980 8679 41180
rect 8759 40980 8789 41180
rect 8869 40980 8899 41180
rect 8979 40980 9009 41180
rect 9089 40980 9119 41180
rect 9199 40980 9229 41180
rect 9309 40980 9339 41180
rect 9419 40980 9449 41180
rect 9529 40980 9559 41180
rect 9639 40980 9669 41180
rect 9749 40980 9779 41180
rect 9859 40980 9889 41180
rect 2719 39760 2749 40560
rect 3049 39760 3079 40560
rect 6419 39660 6449 39860
rect 6529 39660 6559 39860
rect 6639 39660 6669 39860
rect 6749 39660 6779 39860
rect 6859 39660 6889 39860
rect 6969 39660 6999 39860
rect 7079 39660 7109 39860
rect 7189 39660 7219 39860
rect 7299 39660 7329 39860
rect 7409 39660 7439 39860
rect 7519 39660 7549 39860
rect 7629 39660 7659 39860
rect 7739 39660 7769 39860
rect 7849 39660 7879 39860
rect 7959 39660 7989 39860
rect 8069 39660 8099 39860
rect 8179 39660 8209 39860
rect 8289 39660 8319 39860
rect 8399 39660 8429 39860
rect 8509 39660 8539 39860
rect 8619 39660 8649 39860
rect 8729 39660 8759 39860
rect 8839 39660 8869 39860
rect 8949 39660 8979 39860
rect 9059 39660 9089 39860
rect 9169 39660 9199 39860
rect 9279 39660 9309 39860
rect 9389 39660 9419 39860
rect 9499 39660 9529 39860
rect 9609 39660 9639 39860
rect 9719 39660 9749 39860
rect 9829 39660 9859 39860
rect 3840 36250 3870 37050
rect 3950 36250 3980 37050
rect 4060 36250 4090 37050
rect 4170 36250 4200 37050
rect 4280 36250 4310 37050
rect 4390 36250 4420 37050
rect 4650 36250 4680 37050
rect 4760 36250 4790 37050
rect 4870 36250 4900 37050
rect 4980 36250 5010 37050
rect 5090 36250 5120 37050
rect 5200 36250 5230 37050
rect 5530 36650 5560 37050
rect 5640 36650 5670 37050
rect 5750 36650 5780 37050
rect 5860 36650 5890 37050
rect 5970 36650 6000 37050
rect 6080 36650 6110 37050
rect 6410 36390 6440 36590
rect 6520 36390 6550 36590
rect 6770 36190 6800 36590
rect 6880 36190 6910 36590
rect 7030 36190 7060 36590
rect 7140 36190 7170 36590
rect 7370 36390 7400 36590
rect 7480 36390 7510 36590
rect 7750 36390 7780 36590
rect 7860 36390 7890 36590
rect 8130 36390 8160 36590
rect 8240 36390 8270 36590
rect 8510 36390 8540 36590
rect 8620 36390 8650 36590
rect 8850 36190 8880 36590
rect 8960 36190 8990 36590
rect 9110 36190 9140 36590
rect 9220 36190 9250 36590
rect 9450 36390 9480 36590
rect 9560 36390 9590 36590
rect 9830 36390 9860 36590
rect 9940 36390 9970 36590
rect 10210 36390 10240 36590
rect 10320 36390 10350 36590
rect 10590 36390 10620 36590
rect 10700 36390 10730 36590
rect 16530 35610 16560 35840
rect 16640 35610 16670 35840
rect 16750 35610 16780 35840
rect 16860 35610 16890 35840
rect 16970 35610 17000 35840
rect 17080 35610 17110 35840
rect 16530 34450 16560 35350
rect 16640 34450 16670 35350
rect 16750 34450 16780 35350
rect 16860 34450 16890 35350
rect 16970 34450 17000 35350
rect 17080 34450 17110 35350
rect 17420 34960 17450 35160
rect 17820 34910 17850 35110
rect 18360 34960 18390 35160
rect 18760 34960 18790 35160
rect 19830 34950 19860 35150
rect 20080 34950 20110 35150
rect 21490 35610 21520 35840
rect 21600 35610 21630 35840
rect 21710 35610 21740 35840
rect 21820 35610 21850 35840
rect 21930 35610 21960 35840
rect 22040 35610 22070 35840
rect 17640 34440 17670 34640
rect 18100 34440 18130 34640
rect 18580 34440 18610 34640
rect 19040 34440 19070 34640
rect 19370 34450 19400 34850
rect 19830 34370 19860 34570
rect 21100 34450 21130 34850
rect 21490 34450 21520 35350
rect 21600 34450 21630 35350
rect 21710 34450 21740 35350
rect 21820 34450 21850 35350
rect 21930 34450 21960 35350
rect 22040 34450 22070 35350
rect 22380 34960 22410 35160
rect 22780 34910 22810 35110
rect 23320 34960 23350 35160
rect 23720 34960 23750 35160
rect 24790 34950 24820 35150
rect 25040 34950 25070 35150
rect 22600 34440 22630 34640
rect 23060 34440 23090 34640
rect 23540 34440 23570 34640
rect 24000 34440 24030 34640
rect 24330 34450 24360 34850
rect 24790 34370 24820 34570
rect 2240 30800 2270 31600
rect 2350 30800 2380 31600
rect 2460 30800 2490 31600
rect 2570 30800 2600 31600
rect 2680 30800 2710 31600
rect 2790 30800 2820 31600
rect 3050 30800 3080 31600
rect 3160 30800 3190 31600
rect 3270 30800 3300 31600
rect 3380 30800 3410 31600
rect 3490 30800 3520 31600
rect 3600 30800 3630 31600
rect 3930 31200 3960 31600
rect 4040 31200 4070 31600
rect 4150 31200 4180 31600
rect 4260 31200 4290 31600
rect 4370 31200 4400 31600
rect 4480 31200 4510 31600
rect 4790 31200 4820 31600
rect 4900 31200 4930 31600
rect 5010 31200 5040 31600
rect 5120 31200 5150 31600
rect 5230 31200 5260 31600
rect 5340 31200 5370 31600
rect 5650 31200 5680 31600
rect 5760 31200 5790 31600
rect 5870 31200 5900 31600
rect 5980 31200 6010 31600
rect 6090 31200 6120 31600
rect 6200 31200 6230 31600
rect 14178 31360 14208 31660
rect 16530 31550 16560 31780
rect 16640 31550 16670 31780
rect 16750 31550 16780 31780
rect 16860 31550 16890 31780
rect 16970 31550 17000 31780
rect 17080 31550 17110 31780
rect 6470 31040 6500 31240
rect 6580 31040 6610 31240
rect 6830 30840 6860 31240
rect 6940 30840 6970 31240
rect 7090 30840 7120 31240
rect 7200 30840 7230 31240
rect 7430 31040 7460 31240
rect 7540 31040 7570 31240
rect 7810 31040 7840 31240
rect 7920 31040 7950 31240
rect 8190 31040 8220 31240
rect 8300 31040 8330 31240
rect 8570 31040 8600 31240
rect 8680 31040 8710 31240
rect 8910 30840 8940 31240
rect 9020 30840 9050 31240
rect 9170 30840 9200 31240
rect 9280 30840 9310 31240
rect 9510 31040 9540 31240
rect 9620 31040 9650 31240
rect 9890 31040 9920 31240
rect 10000 31040 10030 31240
rect 10270 31040 10300 31240
rect 10380 31040 10410 31240
rect 10650 31040 10680 31240
rect 10760 31040 10790 31240
rect 11030 31040 11060 31240
rect 11140 31040 11170 31240
rect 16530 30390 16560 31290
rect 16640 30390 16670 31290
rect 16750 30390 16780 31290
rect 16860 30390 16890 31290
rect 16970 30390 17000 31290
rect 17080 30390 17110 31290
rect 17420 30900 17450 31100
rect 17820 30850 17850 31050
rect 18360 30900 18390 31100
rect 18760 30900 18790 31100
rect 20090 30890 20120 31090
rect 20340 30890 20370 31090
rect 21550 31540 21580 31770
rect 21660 31540 21690 31770
rect 21770 31540 21800 31770
rect 21880 31540 21910 31770
rect 21990 31540 22020 31770
rect 22100 31540 22130 31770
rect 17640 30380 17670 30580
rect 18100 30380 18130 30580
rect 18580 30380 18610 30580
rect 19040 30380 19070 30580
rect 19370 30390 19400 30790
rect 19630 30390 19660 30790
rect 20090 30310 20120 30510
rect 21160 30390 21190 30790
rect 21550 30380 21580 31280
rect 21660 30380 21690 31280
rect 21770 30380 21800 31280
rect 21880 30380 21910 31280
rect 21990 30380 22020 31280
rect 22100 30380 22130 31280
rect 22440 30890 22470 31090
rect 22840 30840 22870 31040
rect 23380 30890 23410 31090
rect 23780 30890 23810 31090
rect 25050 30880 25080 31080
rect 25300 30880 25330 31080
rect 22660 30370 22690 30570
rect 23120 30370 23150 30570
rect 23600 30370 23630 30570
rect 24060 30370 24090 30570
rect 24390 30380 24420 30780
rect 24650 30380 24680 30780
rect 25050 30300 25080 30500
rect 7390 24370 7420 24570
rect 7500 24370 7530 24570
rect 7920 24370 7950 24570
rect 8030 24370 8060 24570
rect 8550 24360 8580 24760
rect 8700 24360 8730 24760
rect 8930 24630 8960 24830
rect 9290 24360 9320 24560
rect 9400 24360 9430 24560
rect 9630 24360 9660 24760
rect 9740 24360 9770 24760
rect 9890 24360 9920 24760
rect 10000 24360 10030 24760
rect 10230 24360 10260 24560
rect 10340 24360 10370 24560
rect 10620 24360 10650 24760
rect 10730 24360 10760 24760
rect 10880 24360 10910 24760
rect 10990 24360 11020 24760
rect 11220 24360 11250 24560
rect 11330 24360 11360 24560
rect 11620 24360 11650 24760
rect 11730 24360 11760 24760
rect 11880 24360 11910 24760
rect 11990 24360 12020 24760
rect 12950 24640 12980 24840
rect 13180 24640 13210 24840
rect 13290 24640 13320 24840
rect 13520 24640 13550 24840
rect 13630 24640 13660 24840
rect 13740 24640 13770 24840
rect 13850 24640 13880 24840
rect 14080 24640 14110 24840
rect 14190 24640 14220 24840
rect 14300 24640 14330 24840
rect 14410 24640 14440 24840
rect 14520 24640 14550 24840
rect 14630 24640 14660 24840
rect 14740 24640 14770 24840
rect 14850 24640 14880 24840
rect 15140 24640 15170 24840
rect 15250 24640 15280 24840
rect 15360 24640 15390 24840
rect 15470 24640 15500 24840
rect 15580 24640 15610 24840
rect 15690 24640 15720 24840
rect 15800 24640 15830 24840
rect 15910 24640 15940 24840
rect 16020 24640 16050 24840
rect 16130 24640 16160 24840
rect 16240 24640 16270 24840
rect 16350 24640 16380 24840
rect 16460 24640 16490 24840
rect 16570 24640 16600 24840
rect 16680 24640 16710 24840
rect 16790 24640 16820 24840
rect 17090 24640 17120 24840
rect 17200 24640 17230 24840
rect 17310 24640 17340 24840
rect 17420 24640 17450 24840
rect 17530 24640 17560 24840
rect 17640 24640 17670 24840
rect 17750 24640 17780 24840
rect 17860 24640 17890 24840
rect 17970 24640 18000 24840
rect 18080 24640 18110 24840
rect 18190 24640 18220 24840
rect 18300 24640 18330 24840
rect 18410 24640 18440 24840
rect 18520 24640 18550 24840
rect 18630 24640 18660 24840
rect 18740 24640 18770 24840
rect 18850 24640 18880 24840
rect 18960 24640 18990 24840
rect 19070 24640 19100 24840
rect 19180 24640 19210 24840
rect 19290 24640 19320 24840
rect 19400 24640 19430 24840
rect 19510 24640 19540 24840
rect 19620 24640 19650 24840
rect 19730 24640 19760 24840
rect 19840 24640 19870 24840
rect 19950 24640 19980 24840
rect 20060 24640 20090 24840
rect 20170 24640 20200 24840
rect 20280 24640 20310 24840
rect 20390 24640 20420 24840
rect 20500 24640 20530 24840
rect 12220 24360 12250 24560
rect 12330 24360 12360 24560
rect 12600 24360 12630 24560
rect 12710 24360 12740 24560
rect 7430 22810 7460 23210
rect 7540 22810 7570 23210
rect 7690 22810 7720 23210
rect 7800 22810 7830 23210
rect 8030 23010 8060 23210
rect 8140 23010 8170 23210
rect 8550 22810 8580 23210
rect 8700 22810 8730 23210
rect 9290 23010 9320 23210
rect 9400 23010 9430 23210
rect 8930 22740 8960 22940
rect 9630 22810 9660 23210
rect 9740 22810 9770 23210
rect 9890 22810 9920 23210
rect 10000 22810 10030 23210
rect 10230 23010 10260 23210
rect 10340 23010 10370 23210
rect 10620 22810 10650 23210
rect 10730 22810 10760 23210
rect 10880 22810 10910 23210
rect 10990 22810 11020 23210
rect 11220 23010 11250 23210
rect 11330 23010 11360 23210
rect 11620 22810 11650 23210
rect 11730 22810 11760 23210
rect 11880 22810 11910 23210
rect 11990 22810 12020 23210
rect 12220 23010 12250 23210
rect 12330 23010 12360 23210
rect 12600 23010 12630 23210
rect 12710 23010 12740 23210
rect 12950 22730 12980 22930
rect 13180 22730 13210 22930
rect 13290 22730 13320 22930
rect 13520 22730 13550 22930
rect 13630 22730 13660 22930
rect 13740 22730 13770 22930
rect 13850 22730 13880 22930
rect 14080 22730 14110 22930
rect 14190 22730 14220 22930
rect 14300 22730 14330 22930
rect 14410 22730 14440 22930
rect 14520 22730 14550 22930
rect 14630 22730 14660 22930
rect 14740 22730 14770 22930
rect 14850 22730 14880 22930
rect 15140 22730 15170 22930
rect 15250 22730 15280 22930
rect 15360 22730 15390 22930
rect 15470 22730 15500 22930
rect 15580 22730 15610 22930
rect 15690 22730 15720 22930
rect 15800 22730 15830 22930
rect 15910 22730 15940 22930
rect 16020 22730 16050 22930
rect 16130 22730 16160 22930
rect 16240 22730 16270 22930
rect 16350 22730 16380 22930
rect 16460 22730 16490 22930
rect 16570 22730 16600 22930
rect 16680 22730 16710 22930
rect 16790 22730 16820 22930
rect 17090 22730 17120 22930
rect 17200 22730 17230 22930
rect 17310 22730 17340 22930
rect 17420 22730 17450 22930
rect 17530 22730 17560 22930
rect 17640 22730 17670 22930
rect 17750 22730 17780 22930
rect 17860 22730 17890 22930
rect 17970 22730 18000 22930
rect 18080 22730 18110 22930
rect 18190 22730 18220 22930
rect 18300 22730 18330 22930
rect 18410 22730 18440 22930
rect 18520 22730 18550 22930
rect 18630 22730 18660 22930
rect 18740 22730 18770 22930
rect 18850 22730 18880 22930
rect 18960 22730 18990 22930
rect 19070 22730 19100 22930
rect 19180 22730 19210 22930
rect 19290 22730 19320 22930
rect 19400 22730 19430 22930
rect 19510 22730 19540 22930
rect 19620 22730 19650 22930
rect 19730 22730 19760 22930
rect 19840 22730 19870 22930
rect 19950 22730 19980 22930
rect 20060 22730 20090 22930
rect 20170 22730 20200 22930
rect 20280 22730 20310 22930
rect 20390 22730 20420 22930
rect 20500 22730 20530 22930
rect 7350 17780 7380 17980
rect 7460 17780 7490 17980
rect 7610 17780 7640 17980
rect 7720 17780 7750 17980
rect 8020 17780 8050 17980
rect 8130 17780 8160 17980
rect 8550 17770 8580 18170
rect 8700 17770 8730 18170
rect 8930 18040 8960 18240
rect 9290 17770 9320 17970
rect 9400 17770 9430 17970
rect 9630 17770 9660 18170
rect 9740 17770 9770 18170
rect 9890 17770 9920 18170
rect 10000 17770 10030 18170
rect 10230 17770 10260 17970
rect 10340 17770 10370 17970
rect 10620 17770 10650 18170
rect 10730 17770 10760 18170
rect 10880 17770 10910 18170
rect 10990 17770 11020 18170
rect 11220 17770 11250 17970
rect 11330 17770 11360 17970
rect 11620 17770 11650 18170
rect 11730 17770 11760 18170
rect 11880 17770 11910 18170
rect 11990 17770 12020 18170
rect 12950 18050 12980 18250
rect 13180 18050 13210 18250
rect 13290 18050 13320 18250
rect 13520 18050 13550 18250
rect 13630 18050 13660 18250
rect 13740 18050 13770 18250
rect 13850 18050 13880 18250
rect 14080 18050 14110 18250
rect 14190 18050 14220 18250
rect 14300 18050 14330 18250
rect 14410 18050 14440 18250
rect 14520 18050 14550 18250
rect 14630 18050 14660 18250
rect 14740 18050 14770 18250
rect 14850 18050 14880 18250
rect 15140 18050 15170 18250
rect 15250 18050 15280 18250
rect 15360 18050 15390 18250
rect 15470 18050 15500 18250
rect 15580 18050 15610 18250
rect 15690 18050 15720 18250
rect 15800 18050 15830 18250
rect 15910 18050 15940 18250
rect 16020 18050 16050 18250
rect 16130 18050 16160 18250
rect 16240 18050 16270 18250
rect 16350 18050 16380 18250
rect 16460 18050 16490 18250
rect 16570 18050 16600 18250
rect 16680 18050 16710 18250
rect 16790 18050 16820 18250
rect 17090 18050 17120 18250
rect 17200 18050 17230 18250
rect 17310 18050 17340 18250
rect 17420 18050 17450 18250
rect 17530 18050 17560 18250
rect 17640 18050 17670 18250
rect 17750 18050 17780 18250
rect 17860 18050 17890 18250
rect 17970 18050 18000 18250
rect 18080 18050 18110 18250
rect 18190 18050 18220 18250
rect 18300 18050 18330 18250
rect 18410 18050 18440 18250
rect 18520 18050 18550 18250
rect 18630 18050 18660 18250
rect 18740 18050 18770 18250
rect 18850 18050 18880 18250
rect 18960 18050 18990 18250
rect 19070 18050 19100 18250
rect 19180 18050 19210 18250
rect 19290 18050 19320 18250
rect 19400 18050 19430 18250
rect 19510 18050 19540 18250
rect 19620 18050 19650 18250
rect 19730 18050 19760 18250
rect 19840 18050 19870 18250
rect 19950 18050 19980 18250
rect 20060 18050 20090 18250
rect 20170 18050 20200 18250
rect 20280 18050 20310 18250
rect 20390 18050 20420 18250
rect 20500 18050 20530 18250
rect 12220 17770 12250 17970
rect 12330 17770 12360 17970
rect 12600 17770 12630 17970
rect 12710 17770 12740 17970
rect 9830 15350 9860 15550
rect 9940 15350 9970 15550
rect 10370 15150 10400 15550
rect 10480 15150 10510 15550
rect 10630 15150 10660 15550
rect 10740 15150 10770 15550
rect 10970 15350 11000 15550
rect 11080 15350 11110 15550
rect 11360 15150 11390 15550
rect 11470 15150 11500 15550
rect 11620 15150 11650 15550
rect 11730 15150 11760 15550
rect 11960 15350 11990 15550
rect 12070 15350 12100 15550
rect 12360 15150 12390 15550
rect 12470 15150 12500 15550
rect 12620 15150 12650 15550
rect 12730 15150 12760 15550
rect 12960 15350 12990 15550
rect 13070 15350 13100 15550
rect 13310 15070 13340 15270
rect 13540 15070 13570 15270
rect 13650 15070 13680 15270
rect 13880 15070 13910 15270
rect 13990 15070 14020 15270
rect 14100 15070 14130 15270
rect 14210 15070 14240 15270
rect 14440 15070 14470 15270
rect 14550 15070 14580 15270
rect 14660 15070 14690 15270
rect 14770 15070 14800 15270
rect 14880 15070 14910 15270
rect 14990 15070 15020 15270
rect 15100 15070 15130 15270
rect 15210 15070 15240 15270
rect 15500 15070 15530 15270
rect 15610 15070 15640 15270
rect 15720 15070 15750 15270
rect 15830 15070 15860 15270
rect 15940 15070 15970 15270
rect 16050 15070 16080 15270
rect 16160 15070 16190 15270
rect 16270 15070 16300 15270
rect 16380 15070 16410 15270
rect 16490 15070 16520 15270
rect 16600 15070 16630 15270
rect 16710 15070 16740 15270
rect 16820 15070 16850 15270
rect 16930 15070 16960 15270
rect 17040 15070 17070 15270
rect 17150 15070 17180 15270
rect 17450 15070 17480 15270
rect 17560 15070 17590 15270
rect 17670 15070 17700 15270
rect 17780 15070 17810 15270
rect 17890 15070 17920 15270
rect 18000 15070 18030 15270
rect 18110 15070 18140 15270
rect 18220 15070 18250 15270
rect 18330 15070 18360 15270
rect 18440 15070 18470 15270
rect 18550 15070 18580 15270
rect 18660 15070 18690 15270
rect 18770 15070 18800 15270
rect 18880 15070 18910 15270
rect 18990 15070 19020 15270
rect 19100 15070 19130 15270
rect 19210 15070 19240 15270
rect 19320 15070 19350 15270
rect 19430 15070 19460 15270
rect 19540 15070 19570 15270
rect 19650 15070 19680 15270
rect 19760 15070 19790 15270
rect 19870 15070 19900 15270
rect 19980 15070 20010 15270
rect 20090 15070 20120 15270
rect 20200 15070 20230 15270
rect 20310 15070 20340 15270
rect 20420 15070 20450 15270
rect 20530 15070 20560 15270
rect 20640 15070 20670 15270
rect 20750 15070 20780 15270
rect 20860 15070 20890 15270
rect 7350 12120 7380 12320
rect 7460 12120 7490 12320
rect 7870 12120 7900 12520
rect 7980 12120 8010 12520
rect 8130 12120 8160 12520
rect 8240 12120 8270 12520
rect 8620 12080 8650 12480
rect 8770 12080 8800 12480
rect 9000 12390 9030 12590
rect 9260 12390 9290 12590
rect 9510 12390 9540 12590
rect 9930 12120 9960 12320
rect 10040 12120 10070 12320
rect 10470 12120 10500 12520
rect 10580 12120 10610 12520
rect 10730 12120 10760 12520
rect 10840 12120 10870 12520
rect 11070 12120 11100 12320
rect 11180 12120 11210 12320
rect 11460 12120 11490 12520
rect 11570 12120 11600 12520
rect 11720 12120 11750 12520
rect 11830 12120 11860 12520
rect 12060 12120 12090 12320
rect 12170 12120 12200 12320
rect 12460 12120 12490 12520
rect 12570 12120 12600 12520
rect 12720 12120 12750 12520
rect 12830 12120 12860 12520
rect 13410 12400 13440 12600
rect 13640 12400 13670 12600
rect 13750 12400 13780 12600
rect 13980 12400 14010 12600
rect 14090 12400 14120 12600
rect 14200 12400 14230 12600
rect 14310 12400 14340 12600
rect 14540 12400 14570 12600
rect 14650 12400 14680 12600
rect 14760 12400 14790 12600
rect 14870 12400 14900 12600
rect 14980 12400 15010 12600
rect 15090 12400 15120 12600
rect 15200 12400 15230 12600
rect 15310 12400 15340 12600
rect 15600 12400 15630 12600
rect 15710 12400 15740 12600
rect 15820 12400 15850 12600
rect 15930 12400 15960 12600
rect 16040 12400 16070 12600
rect 16150 12400 16180 12600
rect 16260 12400 16290 12600
rect 16370 12400 16400 12600
rect 16480 12400 16510 12600
rect 16590 12400 16620 12600
rect 16700 12400 16730 12600
rect 16810 12400 16840 12600
rect 16920 12400 16950 12600
rect 17030 12400 17060 12600
rect 17140 12400 17170 12600
rect 17250 12400 17280 12600
rect 17550 12400 17580 12600
rect 17660 12400 17690 12600
rect 17770 12400 17800 12600
rect 17880 12400 17910 12600
rect 17990 12400 18020 12600
rect 18100 12400 18130 12600
rect 18210 12400 18240 12600
rect 18320 12400 18350 12600
rect 18430 12400 18460 12600
rect 18540 12400 18570 12600
rect 18650 12400 18680 12600
rect 18760 12400 18790 12600
rect 18870 12400 18900 12600
rect 18980 12400 19010 12600
rect 19090 12400 19120 12600
rect 19200 12400 19230 12600
rect 19310 12400 19340 12600
rect 19420 12400 19450 12600
rect 19530 12400 19560 12600
rect 19640 12400 19670 12600
rect 19750 12400 19780 12600
rect 19860 12400 19890 12600
rect 19970 12400 20000 12600
rect 20080 12400 20110 12600
rect 20190 12400 20220 12600
rect 20300 12400 20330 12600
rect 20410 12400 20440 12600
rect 20520 12400 20550 12600
rect 20630 12400 20660 12600
rect 20740 12400 20770 12600
rect 20850 12400 20880 12600
rect 20960 12400 20990 12600
rect 13060 12120 13090 12320
rect 13170 12120 13200 12320
rect 7920 11100 7950 11300
rect 8030 11100 8060 11300
rect 8180 11100 8210 11300
rect 8290 11100 8320 11300
rect 7350 10730 7380 10930
rect 7460 10730 7490 10930
rect 8710 10580 8740 10980
rect 8860 10580 8890 10980
rect 9930 10730 9960 10930
rect 10040 10730 10070 10930
rect 9090 10470 9120 10670
rect 9350 10470 9380 10670
rect 9600 10470 9630 10670
rect 10470 10530 10500 10930
rect 10580 10530 10610 10930
rect 10730 10530 10760 10930
rect 10840 10530 10870 10930
rect 11070 10730 11100 10930
rect 11180 10730 11210 10930
rect 11460 10530 11490 10930
rect 11570 10530 11600 10930
rect 11720 10530 11750 10930
rect 11830 10530 11860 10930
rect 12060 10730 12090 10930
rect 12170 10730 12200 10930
rect 12460 10530 12490 10930
rect 12570 10530 12600 10930
rect 12720 10530 12750 10930
rect 12830 10530 12860 10930
rect 13060 10730 13090 10930
rect 13170 10730 13200 10930
rect 13400 10450 13430 10650
rect 13630 10450 13660 10650
rect 13740 10450 13770 10650
rect 13970 10450 14000 10650
rect 14080 10450 14110 10650
rect 14190 10450 14220 10650
rect 14300 10450 14330 10650
rect 14530 10450 14560 10650
rect 14640 10450 14670 10650
rect 14750 10450 14780 10650
rect 14860 10450 14890 10650
rect 14970 10450 15000 10650
rect 15080 10450 15110 10650
rect 15190 10450 15220 10650
rect 15300 10450 15330 10650
rect 15590 10450 15620 10650
rect 15700 10450 15730 10650
rect 15810 10450 15840 10650
rect 15920 10450 15950 10650
rect 16030 10450 16060 10650
rect 16140 10450 16170 10650
rect 16250 10450 16280 10650
rect 16360 10450 16390 10650
rect 16470 10450 16500 10650
rect 16580 10450 16610 10650
rect 16690 10450 16720 10650
rect 16800 10450 16830 10650
rect 16910 10450 16940 10650
rect 17020 10450 17050 10650
rect 17130 10450 17160 10650
rect 17240 10450 17270 10650
rect 17540 10450 17570 10650
rect 17650 10450 17680 10650
rect 17760 10450 17790 10650
rect 17870 10450 17900 10650
rect 17980 10450 18010 10650
rect 18090 10450 18120 10650
rect 18200 10450 18230 10650
rect 18310 10450 18340 10650
rect 18420 10450 18450 10650
rect 18530 10450 18560 10650
rect 18640 10450 18670 10650
rect 18750 10450 18780 10650
rect 18860 10450 18890 10650
rect 18970 10450 19000 10650
rect 19080 10450 19110 10650
rect 19190 10450 19220 10650
rect 19300 10450 19330 10650
rect 19410 10450 19440 10650
rect 19520 10450 19550 10650
rect 19630 10450 19660 10650
rect 19740 10450 19770 10650
rect 19850 10450 19880 10650
rect 19960 10450 19990 10650
rect 20070 10450 20100 10650
rect 20180 10450 20210 10650
rect 20290 10450 20320 10650
rect 20400 10450 20430 10650
rect 20510 10450 20540 10650
rect 20620 10450 20650 10650
rect 20730 10450 20760 10650
rect 20840 10450 20870 10650
rect 20950 10450 20980 10650
rect 9940 3210 9970 3810
rect 10050 3210 10080 3810
rect 10160 3210 10190 3810
rect 10270 3210 10300 3810
rect 10380 3210 10410 3810
rect 10490 3210 10520 3810
rect 10600 3210 10630 3810
rect 10710 3210 10740 3810
rect 10820 3210 10850 3810
rect 10930 3210 10960 3810
rect 11040 3210 11070 3810
rect 11150 3210 11180 3810
rect 11260 3210 11290 3810
rect 11370 3210 11400 3810
rect 11480 3210 11510 3810
rect 11590 3210 11620 3810
rect 11700 3210 11730 3810
rect 11810 3210 11840 3810
rect 11920 3210 11950 3810
rect 12030 3210 12060 3810
rect 12140 3210 12170 3810
rect 12250 3210 12280 3810
rect 12360 3210 12390 3810
rect 12470 3210 12500 3810
rect 12580 3210 12610 3810
rect 12690 3210 12720 3810
rect 12800 3210 12830 3810
rect 12910 3210 12940 3810
rect 13020 3210 13050 3810
rect 13130 3210 13160 3810
rect 13700 3540 13730 4140
rect 13810 3540 13840 4140
rect 13920 3540 13950 4140
rect 14030 3540 14060 4140
rect 14140 3540 14170 4140
rect 14250 3540 14280 4140
rect 14360 3540 14390 4140
rect 14470 3540 14500 4140
rect 14580 3540 14610 4140
rect 14690 3540 14720 4140
rect 14800 3540 14830 4140
rect 14910 3540 14940 4140
rect 15020 3540 15050 4140
rect 15130 3540 15160 4140
rect 15240 3540 15270 4140
rect 15350 3540 15380 4140
rect 15460 3540 15490 4140
rect 15570 3540 15600 4140
rect 15680 3540 15710 4140
rect 15790 3540 15820 4140
rect 15900 3540 15930 4140
rect 16010 3540 16040 4140
rect 16120 3540 16150 4140
rect 16230 3540 16260 4140
rect 16340 3540 16370 4140
rect 16450 3540 16480 4140
rect 16560 3540 16590 4140
rect 16670 3540 16700 4140
rect 16780 3540 16810 4140
rect 16890 3540 16920 4140
rect 24350 2670 25350 2700
rect 24350 2560 25350 2590
rect 24350 2450 25350 2480
rect 24350 2340 25350 2370
rect 24350 2230 25350 2260
rect 24350 2120 25350 2150
rect 9960 730 9990 1330
rect 10070 730 10100 1330
rect 10180 730 10210 1330
rect 10290 730 10320 1330
rect 10400 730 10430 1330
rect 10510 730 10540 1330
rect 10620 730 10650 1330
rect 10730 730 10760 1330
rect 10840 730 10870 1330
rect 10950 730 10980 1330
rect 11060 730 11090 1330
rect 11170 730 11200 1330
rect 11280 730 11310 1330
rect 11390 730 11420 1330
rect 11500 730 11530 1330
rect 11610 730 11640 1330
rect 11720 730 11750 1330
rect 11830 730 11860 1330
rect 11940 730 11970 1330
rect 12050 730 12080 1330
rect 12160 730 12190 1330
rect 12270 730 12300 1330
rect 12380 730 12410 1330
rect 12490 730 12520 1330
rect 12600 730 12630 1330
rect 12710 730 12740 1330
rect 12820 730 12850 1330
rect 12930 730 12960 1330
rect 13040 730 13070 1330
rect 13150 730 13180 1330
rect 13700 720 13730 1320
rect 13810 720 13840 1320
rect 13920 720 13950 1320
rect 14030 720 14060 1320
rect 14140 720 14170 1320
rect 14250 720 14280 1320
rect 14360 720 14390 1320
rect 14470 720 14500 1320
rect 14580 720 14610 1320
rect 14690 720 14720 1320
rect 14800 720 14830 1320
rect 14910 720 14940 1320
rect 15020 720 15050 1320
rect 15130 720 15160 1320
rect 15240 720 15270 1320
rect 15350 720 15380 1320
rect 15460 720 15490 1320
rect 15570 720 15600 1320
rect 15680 720 15710 1320
rect 15790 720 15820 1320
rect 15900 720 15930 1320
rect 16010 720 16040 1320
rect 16120 720 16150 1320
rect 16230 720 16260 1320
rect 16340 720 16370 1320
rect 16450 720 16480 1320
rect 16560 720 16590 1320
rect 16670 720 16700 1320
rect 16780 720 16810 1320
rect 16890 720 16920 1320
<< pmos >>
rect 21790 42180 21820 42880
rect 22020 42180 22050 42880
rect 22650 42190 22680 42890
rect 22950 42190 22980 42890
rect 23060 42190 23090 42890
rect 23530 42480 23560 43180
rect 2629 41720 2659 41920
rect 2739 41720 2769 41920
rect 2849 41720 2879 41920
rect 2509 41000 2539 41400
rect 2619 41000 2649 41400
rect 2729 41000 2759 41400
rect 2839 41000 2869 41400
rect 2949 41000 2979 41400
rect 3459 41070 3489 41820
rect 3569 41070 3599 41820
rect 3679 41070 3709 41820
rect 3789 41070 3819 41820
rect 3899 41070 3929 41820
rect 4009 41070 4039 41820
rect 4119 41070 4149 41820
rect 4229 41070 4259 41820
rect 4609 41060 4639 41810
rect 4719 41060 4749 41810
rect 4829 41060 4859 41810
rect 4939 41060 4969 41810
rect 5049 41060 5079 41810
rect 5159 41060 5189 41810
rect 5269 41060 5299 41810
rect 5379 41060 5409 41810
rect 6019 41340 6049 41840
rect 6249 41340 6279 41840
rect 6359 41340 6389 41840
rect 6589 41340 6619 41840
rect 6699 41340 6729 41840
rect 6809 41340 6839 41840
rect 6919 41340 6949 41840
rect 7149 41340 7179 41840
rect 7259 41340 7289 41840
rect 7369 41340 7399 41840
rect 7479 41340 7509 41840
rect 7589 41340 7619 41840
rect 7699 41340 7729 41840
rect 7809 41340 7839 41840
rect 7919 41340 7949 41840
rect 8209 41340 8239 41840
rect 8319 41340 8349 41840
rect 8429 41340 8459 41840
rect 8539 41340 8569 41840
rect 8649 41340 8679 41840
rect 8759 41340 8789 41840
rect 8869 41340 8899 41840
rect 8979 41340 9009 41840
rect 9089 41340 9119 41840
rect 9199 41340 9229 41840
rect 9309 41340 9339 41840
rect 9419 41340 9449 41840
rect 9529 41340 9559 41840
rect 9639 41340 9669 41840
rect 9749 41340 9779 41840
rect 9859 41340 9889 41840
rect 3329 39780 3359 40530
rect 3439 39780 3469 40530
rect 3549 39780 3579 40530
rect 3659 39780 3689 40530
rect 3769 39780 3799 40530
rect 3879 39780 3909 40530
rect 3989 39780 4019 40530
rect 4099 39780 4129 40530
rect 4609 39780 4639 40530
rect 4719 39780 4749 40530
rect 4829 39780 4859 40530
rect 4939 39780 4969 40530
rect 5049 39780 5079 40530
rect 5159 39780 5189 40530
rect 5269 39780 5299 40530
rect 5379 39780 5409 40530
rect 6419 40020 6449 40520
rect 6529 40020 6559 40520
rect 6639 40020 6669 40520
rect 6749 40020 6779 40520
rect 6859 40020 6889 40520
rect 6969 40020 6999 40520
rect 7079 40020 7109 40520
rect 7189 40020 7219 40520
rect 7299 40020 7329 40520
rect 7409 40020 7439 40520
rect 7519 40020 7549 40520
rect 7629 40020 7659 40520
rect 7739 40020 7769 40520
rect 7849 40020 7879 40520
rect 7959 40020 7989 40520
rect 8069 40020 8099 40520
rect 8179 40020 8209 40520
rect 8289 40020 8319 40520
rect 8399 40020 8429 40520
rect 8509 40020 8539 40520
rect 8619 40020 8649 40520
rect 8729 40020 8759 40520
rect 8839 40020 8869 40520
rect 8949 40020 8979 40520
rect 9059 40020 9089 40520
rect 9169 40020 9199 40520
rect 9279 40020 9309 40520
rect 9389 40020 9419 40520
rect 9499 40020 9529 40520
rect 9609 40020 9639 40520
rect 9719 40020 9749 40520
rect 9829 40020 9859 40520
rect 3840 33690 3870 34690
rect 3950 33690 3980 34690
rect 4060 33690 4090 34690
rect 4170 33690 4200 34690
rect 4280 33690 4310 34690
rect 4390 33690 4420 34690
rect 4650 33690 4680 34690
rect 4760 33690 4790 34690
rect 4870 33690 4900 34690
rect 4980 33690 5010 34690
rect 5090 33690 5120 34690
rect 5200 33690 5230 34690
rect 5530 33760 5560 34760
rect 5640 33760 5670 34760
rect 5750 33760 5780 34760
rect 5860 33760 5890 34760
rect 5970 33760 6000 34760
rect 6080 33760 6110 34760
rect 6410 34260 6440 34760
rect 6520 34260 6550 34760
rect 15410 35770 15440 35970
rect 15520 35770 15550 35970
rect 17530 35580 17560 36080
rect 17780 35580 17810 36080
rect 18100 35580 18130 36080
rect 18470 35580 18500 36080
rect 18720 35580 18750 36080
rect 19040 35580 19070 36080
rect 6770 34250 6800 34750
rect 6880 34250 6910 34750
rect 7030 34250 7060 34750
rect 7140 34250 7170 34750
rect 7370 34250 7400 34750
rect 7480 34250 7510 34750
rect 7750 34250 7780 34750
rect 7860 34250 7890 34750
rect 8130 34250 8160 34750
rect 8240 34250 8270 34750
rect 8510 34250 8540 34750
rect 8620 34250 8650 34750
rect 8850 34250 8880 34750
rect 8960 34250 8990 34750
rect 9110 34250 9140 34750
rect 9220 34250 9250 34750
rect 9450 34250 9480 34750
rect 9560 34250 9590 34750
rect 9830 34250 9860 34750
rect 9940 34250 9970 34750
rect 10210 34250 10240 34750
rect 10320 34250 10350 34750
rect 10590 34250 10620 34750
rect 10700 34250 10730 34750
rect 19370 35010 19400 36010
rect 19830 35600 19860 36100
rect 20080 35600 20110 36100
rect 21100 35010 21130 36010
rect 22490 35580 22520 36080
rect 22740 35580 22770 36080
rect 23060 35580 23090 36080
rect 23430 35580 23460 36080
rect 23680 35580 23710 36080
rect 24000 35580 24030 36080
rect 24330 35010 24360 36010
rect 24790 35600 24820 36100
rect 25040 35600 25070 36100
rect 13958 32040 13988 32240
rect 14068 32040 14098 32240
rect 14178 32040 14208 32240
rect 17530 31520 17560 32020
rect 17780 31520 17810 32020
rect 18100 31520 18130 32020
rect 18470 31520 18500 32020
rect 18720 31520 18750 32020
rect 19040 31520 19070 32020
rect 2240 29440 2270 30440
rect 2350 29440 2380 30440
rect 2460 29440 2490 30440
rect 2570 29440 2600 30440
rect 2680 29440 2710 30440
rect 2790 29440 2820 30440
rect 3050 29440 3080 30440
rect 3160 29440 3190 30440
rect 3270 29440 3300 30440
rect 3380 29440 3410 30440
rect 3490 29440 3520 30440
rect 3600 29440 3630 30440
rect 3930 29510 3960 30510
rect 4040 29510 4070 30510
rect 4150 29510 4180 30510
rect 4260 29510 4290 30510
rect 4370 29510 4400 30510
rect 4480 29510 4510 30510
rect 4790 29510 4820 30510
rect 4900 29510 4930 30510
rect 5010 29510 5040 30510
rect 5120 29510 5150 30510
rect 5230 29510 5260 30510
rect 5340 29510 5370 30510
rect 5650 29510 5680 30510
rect 5760 29510 5790 30510
rect 5870 29510 5900 30510
rect 5980 29510 6010 30510
rect 6090 29510 6120 30510
rect 6200 29510 6230 30510
rect 6470 30110 6500 30610
rect 6580 30110 6610 30610
rect 6830 30100 6860 30600
rect 6940 30100 6970 30600
rect 7090 30100 7120 30600
rect 7200 30100 7230 30600
rect 7430 30100 7460 30600
rect 7540 30100 7570 30600
rect 7810 30100 7840 30600
rect 7920 30100 7950 30600
rect 8190 30100 8220 30600
rect 8300 30100 8330 30600
rect 8570 30100 8600 30600
rect 8680 30100 8710 30600
rect 8910 30100 8940 30600
rect 9020 30100 9050 30600
rect 9170 30100 9200 30600
rect 9280 30100 9310 30600
rect 9510 30100 9540 30600
rect 9620 30100 9650 30600
rect 9890 30100 9920 30600
rect 10000 30100 10030 30600
rect 10270 30100 10300 30600
rect 10380 30100 10410 30600
rect 10650 30100 10680 30600
rect 10760 30100 10790 30600
rect 11030 30100 11060 30600
rect 11140 30100 11170 30600
rect 19370 30950 19400 31950
rect 19630 30950 19660 31950
rect 20090 31520 20120 32020
rect 20340 31520 20370 32020
rect 21160 30950 21190 31950
rect 22550 31510 22580 32010
rect 22800 31510 22830 32010
rect 23120 31510 23150 32010
rect 23490 31510 23520 32010
rect 23740 31510 23770 32010
rect 24060 31510 24090 32010
rect 24390 30940 24420 31940
rect 24650 30940 24680 31940
rect 25050 31530 25080 32030
rect 25300 31530 25330 32030
rect 7390 25990 7420 26490
rect 7500 25990 7530 26490
rect 7920 25990 7950 26490
rect 8030 25990 8060 26490
rect 8550 26000 8580 26500
rect 8700 26000 8730 26500
rect 8930 26000 8960 26500
rect 9290 26000 9320 26500
rect 9400 26000 9430 26500
rect 9630 26000 9660 26500
rect 9740 26000 9770 26500
rect 9890 26000 9920 26500
rect 10000 26000 10030 26500
rect 10230 26000 10260 26500
rect 10340 26000 10370 26500
rect 10620 26000 10650 26500
rect 10730 26000 10760 26500
rect 10880 26000 10910 26500
rect 10990 26000 11020 26500
rect 11220 26000 11250 26500
rect 11330 26000 11360 26500
rect 11620 26000 11650 26500
rect 11730 26000 11760 26500
rect 11880 26000 11910 26500
rect 11990 26000 12020 26500
rect 12220 26000 12250 26500
rect 12330 26000 12360 26500
rect 12600 26000 12630 26500
rect 12710 26000 12740 26500
rect 12950 26000 12980 26500
rect 13180 26000 13210 26500
rect 13290 26000 13320 26500
rect 13520 26000 13550 26500
rect 13630 26000 13660 26500
rect 13740 26000 13770 26500
rect 13850 26000 13880 26500
rect 14080 26000 14110 26500
rect 14190 26000 14220 26500
rect 14300 26000 14330 26500
rect 14410 26000 14440 26500
rect 14520 26000 14550 26500
rect 14630 26000 14660 26500
rect 14740 26000 14770 26500
rect 14850 26000 14880 26500
rect 15140 26000 15170 26500
rect 15250 26000 15280 26500
rect 15360 26000 15390 26500
rect 15470 26000 15500 26500
rect 15580 26000 15610 26500
rect 15690 26000 15720 26500
rect 15800 26000 15830 26500
rect 15910 26000 15940 26500
rect 16020 26000 16050 26500
rect 16130 26000 16160 26500
rect 16240 26000 16270 26500
rect 16350 26000 16380 26500
rect 16460 26000 16490 26500
rect 16570 26000 16600 26500
rect 16680 26000 16710 26500
rect 16790 26000 16820 26500
rect 17090 26000 17120 26500
rect 17200 26000 17230 26500
rect 17310 26000 17340 26500
rect 17420 26000 17450 26500
rect 17530 26000 17560 26500
rect 17640 26000 17670 26500
rect 17750 26000 17780 26500
rect 17860 26000 17890 26500
rect 17970 26000 18000 26500
rect 18080 26000 18110 26500
rect 18190 26000 18220 26500
rect 18300 26000 18330 26500
rect 18410 26000 18440 26500
rect 18520 26000 18550 26500
rect 18630 26000 18660 26500
rect 18740 26000 18770 26500
rect 18850 26000 18880 26500
rect 18960 26000 18990 26500
rect 19070 26000 19100 26500
rect 19180 26000 19210 26500
rect 19290 26000 19320 26500
rect 19400 26000 19430 26500
rect 19510 26000 19540 26500
rect 19620 26000 19650 26500
rect 19730 26000 19760 26500
rect 19840 26000 19870 26500
rect 19950 26000 19980 26500
rect 20060 26000 20090 26500
rect 20170 26000 20200 26500
rect 20280 26000 20310 26500
rect 20390 26000 20420 26500
rect 20500 26000 20530 26500
rect 7430 21080 7460 21580
rect 7540 21080 7570 21580
rect 7690 21080 7720 21580
rect 7800 21080 7830 21580
rect 8030 21080 8060 21580
rect 8140 21080 8170 21580
rect 8550 21070 8580 21570
rect 8700 21070 8730 21570
rect 8930 21070 8960 21570
rect 9290 21070 9320 21570
rect 9400 21070 9430 21570
rect 9630 21070 9660 21570
rect 9740 21070 9770 21570
rect 9890 21070 9920 21570
rect 10000 21070 10030 21570
rect 10230 21070 10260 21570
rect 10340 21070 10370 21570
rect 10620 21070 10650 21570
rect 10730 21070 10760 21570
rect 10880 21070 10910 21570
rect 10990 21070 11020 21570
rect 11220 21070 11250 21570
rect 11330 21070 11360 21570
rect 11620 21070 11650 21570
rect 11730 21070 11760 21570
rect 11880 21070 11910 21570
rect 11990 21070 12020 21570
rect 12220 21070 12250 21570
rect 12330 21070 12360 21570
rect 12600 21070 12630 21570
rect 12710 21070 12740 21570
rect 12950 21070 12980 21570
rect 13180 21070 13210 21570
rect 13290 21070 13320 21570
rect 13520 21070 13550 21570
rect 13630 21070 13660 21570
rect 13740 21070 13770 21570
rect 13850 21070 13880 21570
rect 14080 21070 14110 21570
rect 14190 21070 14220 21570
rect 14300 21070 14330 21570
rect 14410 21070 14440 21570
rect 14520 21070 14550 21570
rect 14630 21070 14660 21570
rect 14740 21070 14770 21570
rect 14850 21070 14880 21570
rect 15140 21070 15170 21570
rect 15250 21070 15280 21570
rect 15360 21070 15390 21570
rect 15470 21070 15500 21570
rect 15580 21070 15610 21570
rect 15690 21070 15720 21570
rect 15800 21070 15830 21570
rect 15910 21070 15940 21570
rect 16020 21070 16050 21570
rect 16130 21070 16160 21570
rect 16240 21070 16270 21570
rect 16350 21070 16380 21570
rect 16460 21070 16490 21570
rect 16570 21070 16600 21570
rect 16680 21070 16710 21570
rect 16790 21070 16820 21570
rect 17090 21070 17120 21570
rect 17200 21070 17230 21570
rect 17310 21070 17340 21570
rect 17420 21070 17450 21570
rect 17530 21070 17560 21570
rect 17640 21070 17670 21570
rect 17750 21070 17780 21570
rect 17860 21070 17890 21570
rect 17970 21070 18000 21570
rect 18080 21070 18110 21570
rect 18190 21070 18220 21570
rect 18300 21070 18330 21570
rect 18410 21070 18440 21570
rect 18520 21070 18550 21570
rect 18630 21070 18660 21570
rect 18740 21070 18770 21570
rect 18850 21070 18880 21570
rect 18960 21070 18990 21570
rect 19070 21070 19100 21570
rect 19180 21070 19210 21570
rect 19290 21070 19320 21570
rect 19400 21070 19430 21570
rect 19510 21070 19540 21570
rect 19620 21070 19650 21570
rect 19730 21070 19760 21570
rect 19840 21070 19870 21570
rect 19950 21070 19980 21570
rect 20060 21070 20090 21570
rect 20170 21070 20200 21570
rect 20280 21070 20310 21570
rect 20390 21070 20420 21570
rect 20500 21070 20530 21570
rect 7350 19360 7380 20360
rect 7460 19360 7490 20360
rect 7610 19360 7640 20360
rect 7720 19360 7750 20360
rect 8020 19860 8050 20360
rect 8130 19860 8160 20360
rect 8550 19410 8580 19910
rect 8700 19410 8730 19910
rect 8930 19410 8960 19910
rect 9290 19410 9320 19910
rect 9400 19410 9430 19910
rect 9630 19410 9660 19910
rect 9740 19410 9770 19910
rect 9890 19410 9920 19910
rect 10000 19410 10030 19910
rect 10230 19410 10260 19910
rect 10340 19410 10370 19910
rect 10620 19410 10650 19910
rect 10730 19410 10760 19910
rect 10880 19410 10910 19910
rect 10990 19410 11020 19910
rect 11220 19410 11250 19910
rect 11330 19410 11360 19910
rect 11620 19410 11650 19910
rect 11730 19410 11760 19910
rect 11880 19410 11910 19910
rect 11990 19410 12020 19910
rect 12220 19410 12250 19910
rect 12330 19410 12360 19910
rect 12600 19410 12630 19910
rect 12710 19410 12740 19910
rect 12950 19410 12980 19910
rect 13180 19410 13210 19910
rect 13290 19410 13320 19910
rect 13520 19410 13550 19910
rect 13630 19410 13660 19910
rect 13740 19410 13770 19910
rect 13850 19410 13880 19910
rect 14080 19410 14110 19910
rect 14190 19410 14220 19910
rect 14300 19410 14330 19910
rect 14410 19410 14440 19910
rect 14520 19410 14550 19910
rect 14630 19410 14660 19910
rect 14740 19410 14770 19910
rect 14850 19410 14880 19910
rect 15140 19410 15170 19910
rect 15250 19410 15280 19910
rect 15360 19410 15390 19910
rect 15470 19410 15500 19910
rect 15580 19410 15610 19910
rect 15690 19410 15720 19910
rect 15800 19410 15830 19910
rect 15910 19410 15940 19910
rect 16020 19410 16050 19910
rect 16130 19410 16160 19910
rect 16240 19410 16270 19910
rect 16350 19410 16380 19910
rect 16460 19410 16490 19910
rect 16570 19410 16600 19910
rect 16680 19410 16710 19910
rect 16790 19410 16820 19910
rect 17090 19410 17120 19910
rect 17200 19410 17230 19910
rect 17310 19410 17340 19910
rect 17420 19410 17450 19910
rect 17530 19410 17560 19910
rect 17640 19410 17670 19910
rect 17750 19410 17780 19910
rect 17860 19410 17890 19910
rect 17970 19410 18000 19910
rect 18080 19410 18110 19910
rect 18190 19410 18220 19910
rect 18300 19410 18330 19910
rect 18410 19410 18440 19910
rect 18520 19410 18550 19910
rect 18630 19410 18660 19910
rect 18740 19410 18770 19910
rect 18850 19410 18880 19910
rect 18960 19410 18990 19910
rect 19070 19410 19100 19910
rect 19180 19410 19210 19910
rect 19290 19410 19320 19910
rect 19400 19410 19430 19910
rect 19510 19410 19540 19910
rect 19620 19410 19650 19910
rect 19730 19410 19760 19910
rect 19840 19410 19870 19910
rect 19950 19410 19980 19910
rect 20060 19410 20090 19910
rect 20170 19410 20200 19910
rect 20280 19410 20310 19910
rect 20390 19410 20420 19910
rect 20500 19410 20530 19910
rect 9830 14410 9860 14910
rect 9940 14410 9970 14910
rect 10370 14410 10400 14910
rect 10480 14410 10510 14910
rect 10630 14410 10660 14910
rect 10740 14410 10770 14910
rect 10970 14410 11000 14910
rect 11080 14410 11110 14910
rect 11360 14410 11390 14910
rect 11470 14410 11500 14910
rect 11620 14410 11650 14910
rect 11730 14410 11760 14910
rect 11960 14410 11990 14910
rect 12070 14410 12100 14910
rect 12360 14410 12390 14910
rect 12470 14410 12500 14910
rect 12620 14410 12650 14910
rect 12730 14410 12760 14910
rect 12960 14410 12990 14910
rect 13070 14410 13100 14910
rect 13310 14410 13340 14910
rect 13540 14410 13570 14910
rect 13650 14410 13680 14910
rect 13880 14410 13910 14910
rect 13990 14410 14020 14910
rect 14100 14410 14130 14910
rect 14210 14410 14240 14910
rect 14440 14410 14470 14910
rect 14550 14410 14580 14910
rect 14660 14410 14690 14910
rect 14770 14410 14800 14910
rect 14880 14410 14910 14910
rect 14990 14410 15020 14910
rect 15100 14410 15130 14910
rect 15210 14410 15240 14910
rect 15500 14410 15530 14910
rect 15610 14410 15640 14910
rect 15720 14410 15750 14910
rect 15830 14410 15860 14910
rect 15940 14410 15970 14910
rect 16050 14410 16080 14910
rect 16160 14410 16190 14910
rect 16270 14410 16300 14910
rect 16380 14410 16410 14910
rect 16490 14410 16520 14910
rect 16600 14410 16630 14910
rect 16710 14410 16740 14910
rect 16820 14410 16850 14910
rect 16930 14410 16960 14910
rect 17040 14410 17070 14910
rect 17150 14410 17180 14910
rect 17450 14410 17480 14910
rect 17560 14410 17590 14910
rect 17670 14410 17700 14910
rect 17780 14410 17810 14910
rect 17890 14410 17920 14910
rect 18000 14410 18030 14910
rect 18110 14410 18140 14910
rect 18220 14410 18250 14910
rect 18330 14410 18360 14910
rect 18440 14410 18470 14910
rect 18550 14410 18580 14910
rect 18660 14410 18690 14910
rect 18770 14410 18800 14910
rect 18880 14410 18910 14910
rect 18990 14410 19020 14910
rect 19100 14410 19130 14910
rect 19210 14410 19240 14910
rect 19320 14410 19350 14910
rect 19430 14410 19460 14910
rect 19540 14410 19570 14910
rect 19650 14410 19680 14910
rect 19760 14410 19790 14910
rect 19870 14410 19900 14910
rect 19980 14410 20010 14910
rect 20090 14410 20120 14910
rect 20200 14410 20230 14910
rect 20310 14410 20340 14910
rect 20420 14410 20450 14910
rect 20530 14410 20560 14910
rect 20640 14410 20670 14910
rect 20750 14410 20780 14910
rect 20860 14410 20890 14910
rect 7350 12760 7380 13260
rect 7460 12760 7490 13260
rect 7870 12760 7900 13260
rect 7980 12760 8010 13260
rect 8130 12760 8160 13260
rect 8240 12760 8270 13260
rect 8620 12760 8650 13260
rect 8770 12760 8800 13260
rect 9000 12760 9030 13260
rect 9260 12760 9290 13260
rect 9510 12760 9540 13260
rect 9930 12760 9960 13260
rect 10040 12760 10070 13260
rect 10470 12760 10500 13260
rect 10580 12760 10610 13260
rect 10730 12760 10760 13260
rect 10840 12760 10870 13260
rect 11070 12760 11100 13260
rect 11180 12760 11210 13260
rect 11460 12760 11490 13260
rect 11570 12760 11600 13260
rect 11720 12760 11750 13260
rect 11830 12760 11860 13260
rect 12060 12760 12090 13260
rect 12170 12760 12200 13260
rect 12460 12760 12490 13260
rect 12570 12760 12600 13260
rect 12720 12760 12750 13260
rect 12830 12760 12860 13260
rect 13060 12760 13090 13260
rect 13170 12760 13200 13260
rect 13410 12760 13440 13260
rect 13640 12760 13670 13260
rect 13750 12760 13780 13260
rect 13980 12760 14010 13260
rect 14090 12760 14120 13260
rect 14200 12760 14230 13260
rect 14310 12760 14340 13260
rect 14540 12760 14570 13260
rect 14650 12760 14680 13260
rect 14760 12760 14790 13260
rect 14870 12760 14900 13260
rect 14980 12760 15010 13260
rect 15090 12760 15120 13260
rect 15200 12760 15230 13260
rect 15310 12760 15340 13260
rect 15600 12760 15630 13260
rect 15710 12760 15740 13260
rect 15820 12760 15850 13260
rect 15930 12760 15960 13260
rect 16040 12760 16070 13260
rect 16150 12760 16180 13260
rect 16260 12760 16290 13260
rect 16370 12760 16400 13260
rect 16480 12760 16510 13260
rect 16590 12760 16620 13260
rect 16700 12760 16730 13260
rect 16810 12760 16840 13260
rect 16920 12760 16950 13260
rect 17030 12760 17060 13260
rect 17140 12760 17170 13260
rect 17250 12760 17280 13260
rect 17550 12760 17580 13260
rect 17660 12760 17690 13260
rect 17770 12760 17800 13260
rect 17880 12760 17910 13260
rect 17990 12760 18020 13260
rect 18100 12760 18130 13260
rect 18210 12760 18240 13260
rect 18320 12760 18350 13260
rect 18430 12760 18460 13260
rect 18540 12760 18570 13260
rect 18650 12760 18680 13260
rect 18760 12760 18790 13260
rect 18870 12760 18900 13260
rect 18980 12760 19010 13260
rect 19090 12760 19120 13260
rect 19200 12760 19230 13260
rect 19310 12760 19340 13260
rect 19420 12760 19450 13260
rect 19530 12760 19560 13260
rect 19640 12760 19670 13260
rect 19750 12760 19780 13260
rect 19860 12760 19890 13260
rect 19970 12760 20000 13260
rect 20080 12760 20110 13260
rect 20190 12760 20220 13260
rect 20300 12760 20330 13260
rect 20410 12760 20440 13260
rect 20520 12760 20550 13260
rect 20630 12760 20660 13260
rect 20740 12760 20770 13260
rect 20850 12760 20880 13260
rect 20960 12760 20990 13260
rect 7350 9790 7380 10290
rect 7460 9790 7490 10290
rect 7920 9720 7950 10720
rect 8030 9720 8060 10720
rect 8180 9720 8210 10720
rect 8290 9720 8320 10720
rect 8710 9800 8740 10300
rect 8860 9800 8890 10300
rect 9090 9800 9120 10300
rect 9350 9800 9380 10300
rect 9600 9800 9630 10300
rect 9930 9790 9960 10290
rect 10040 9790 10070 10290
rect 10470 9790 10500 10290
rect 10580 9790 10610 10290
rect 10730 9790 10760 10290
rect 10840 9790 10870 10290
rect 11070 9790 11100 10290
rect 11180 9790 11210 10290
rect 11460 9790 11490 10290
rect 11570 9790 11600 10290
rect 11720 9790 11750 10290
rect 11830 9790 11860 10290
rect 12060 9790 12090 10290
rect 12170 9790 12200 10290
rect 12460 9790 12490 10290
rect 12570 9790 12600 10290
rect 12720 9790 12750 10290
rect 12830 9790 12860 10290
rect 13060 9790 13090 10290
rect 13170 9790 13200 10290
rect 13400 9790 13430 10290
rect 13630 9790 13660 10290
rect 13740 9790 13770 10290
rect 13970 9790 14000 10290
rect 14080 9790 14110 10290
rect 14190 9790 14220 10290
rect 14300 9790 14330 10290
rect 14530 9790 14560 10290
rect 14640 9790 14670 10290
rect 14750 9790 14780 10290
rect 14860 9790 14890 10290
rect 14970 9790 15000 10290
rect 15080 9790 15110 10290
rect 15190 9790 15220 10290
rect 15300 9790 15330 10290
rect 15590 9790 15620 10290
rect 15700 9790 15730 10290
rect 15810 9790 15840 10290
rect 15920 9790 15950 10290
rect 16030 9790 16060 10290
rect 16140 9790 16170 10290
rect 16250 9790 16280 10290
rect 16360 9790 16390 10290
rect 16470 9790 16500 10290
rect 16580 9790 16610 10290
rect 16690 9790 16720 10290
rect 16800 9790 16830 10290
rect 16910 9790 16940 10290
rect 17020 9790 17050 10290
rect 17130 9790 17160 10290
rect 17240 9790 17270 10290
rect 17540 9790 17570 10290
rect 17650 9790 17680 10290
rect 17760 9790 17790 10290
rect 17870 9790 17900 10290
rect 17980 9790 18010 10290
rect 18090 9790 18120 10290
rect 18200 9790 18230 10290
rect 18310 9790 18340 10290
rect 18420 9790 18450 10290
rect 18530 9790 18560 10290
rect 18640 9790 18670 10290
rect 18750 9790 18780 10290
rect 18860 9790 18890 10290
rect 18970 9790 19000 10290
rect 19080 9790 19110 10290
rect 19190 9790 19220 10290
rect 19300 9790 19330 10290
rect 19410 9790 19440 10290
rect 19520 9790 19550 10290
rect 19630 9790 19660 10290
rect 19740 9790 19770 10290
rect 19850 9790 19880 10290
rect 19960 9790 19990 10290
rect 20070 9790 20100 10290
rect 20180 9790 20210 10290
rect 20290 9790 20320 10290
rect 20400 9790 20430 10290
rect 20510 9790 20540 10290
rect 20620 9790 20650 10290
rect 20730 9790 20760 10290
rect 20840 9790 20870 10290
rect 20950 9790 20980 10290
rect 9970 7060 10000 8260
rect 10080 7060 10110 8260
rect 10190 7060 10220 8260
rect 10300 7060 10330 8260
rect 10410 7060 10440 8260
rect 10520 7060 10550 8260
rect 10630 7060 10660 8260
rect 10740 7060 10770 8260
rect 10850 7060 10880 8260
rect 10960 7060 10990 8260
rect 11070 7060 11100 8260
rect 11180 7060 11210 8260
rect 11290 7060 11320 8260
rect 11400 7060 11430 8260
rect 11510 7060 11540 8260
rect 11620 7060 11650 8260
rect 11730 7060 11760 8260
rect 11840 7060 11870 8260
rect 11950 7060 11980 8260
rect 12060 7060 12090 8260
rect 12170 7060 12200 8260
rect 12280 7060 12310 8260
rect 12390 7060 12420 8260
rect 12500 7060 12530 8260
rect 12610 7060 12640 8260
rect 12720 7060 12750 8260
rect 12830 7060 12860 8260
rect 12940 7060 12970 8260
rect 13050 7060 13080 8260
rect 13160 7060 13190 8260
rect 13740 7060 13770 8260
rect 13850 7060 13880 8260
rect 13960 7060 13990 8260
rect 14070 7060 14100 8260
rect 14180 7060 14210 8260
rect 14290 7060 14320 8260
rect 14400 7060 14430 8260
rect 14510 7060 14540 8260
rect 14620 7060 14650 8260
rect 14730 7060 14760 8260
rect 14840 7060 14870 8260
rect 14950 7060 14980 8260
rect 15060 7060 15090 8260
rect 15170 7060 15200 8260
rect 15280 7060 15310 8260
rect 15390 7060 15420 8260
rect 15500 7060 15530 8260
rect 15610 7060 15640 8260
rect 15720 7060 15750 8260
rect 15830 7060 15860 8260
rect 15940 7060 15970 8260
rect 16050 7060 16080 8260
rect 16160 7060 16190 8260
rect 16270 7060 16300 8260
rect 16380 7060 16410 8260
rect 16490 7060 16520 8260
rect 16600 7060 16630 8260
rect 16710 7060 16740 8260
rect 16820 7060 16850 8260
rect 16930 7060 16960 8260
rect 9940 4420 9970 5620
rect 10050 4420 10080 5620
rect 10160 4420 10190 5620
rect 10270 4420 10300 5620
rect 10380 4420 10410 5620
rect 10490 4420 10520 5620
rect 10600 4420 10630 5620
rect 10710 4420 10740 5620
rect 10820 4420 10850 5620
rect 10930 4420 10960 5620
rect 11040 4420 11070 5620
rect 11150 4420 11180 5620
rect 11260 4420 11290 5620
rect 11370 4420 11400 5620
rect 11480 4420 11510 5620
rect 11590 4420 11620 5620
rect 11700 4420 11730 5620
rect 11810 4420 11840 5620
rect 11920 4420 11950 5620
rect 12030 4420 12060 5620
rect 12140 4420 12170 5620
rect 12250 4420 12280 5620
rect 12360 4420 12390 5620
rect 12470 4420 12500 5620
rect 12580 4420 12610 5620
rect 12690 4420 12720 5620
rect 12800 4420 12830 5620
rect 12910 4420 12940 5620
rect 13020 4420 13050 5620
rect 13130 4420 13160 5620
rect 13700 4660 13730 5860
rect 13810 4660 13840 5860
rect 13920 4660 13950 5860
rect 14030 4660 14060 5860
rect 14140 4660 14170 5860
rect 14250 4660 14280 5860
rect 14360 4660 14390 5860
rect 14470 4660 14500 5860
rect 14580 4660 14610 5860
rect 14690 4660 14720 5860
rect 14800 4660 14830 5860
rect 14910 4660 14940 5860
rect 15020 4660 15050 5860
rect 15130 4660 15160 5860
rect 15240 4660 15270 5860
rect 15350 4660 15380 5860
rect 15460 4660 15490 5860
rect 15570 4660 15600 5860
rect 15680 4660 15710 5860
rect 15790 4660 15820 5860
rect 15900 4660 15930 5860
rect 16010 4660 16040 5860
rect 16120 4660 16150 5860
rect 16230 4660 16260 5860
rect 16340 4660 16370 5860
rect 16450 4660 16480 5860
rect 16560 4660 16590 5860
rect 16670 4660 16700 5860
rect 16780 4660 16810 5860
rect 16890 4660 16920 5860
<< ndiff >>
rect 23370 42080 23450 42100
rect 23370 41920 23390 42080
rect 23430 41920 23450 42080
rect 21720 41860 21790 41880
rect 21720 41700 21730 41860
rect 21770 41700 21790 41860
rect 21720 41680 21790 41700
rect 21820 41860 21890 41880
rect 21820 41700 21840 41860
rect 21880 41700 21890 41860
rect 23370 41900 23450 41920
rect 23480 42080 23550 42100
rect 23480 41920 23500 42080
rect 23540 41920 23550 42080
rect 23480 41900 23550 41920
rect 21820 41680 21890 41700
rect 22580 41690 22650 41710
rect 22580 41530 22590 41690
rect 22630 41530 22650 41690
rect 22580 41510 22650 41530
rect 22680 41690 22750 41710
rect 22680 41530 22700 41690
rect 22740 41530 22750 41690
rect 22680 41510 22750 41530
rect 22880 41690 22950 41710
rect 22880 41530 22890 41690
rect 22930 41530 22950 41690
rect 22880 41510 22950 41530
rect 22980 41690 23060 41710
rect 22980 41530 23000 41690
rect 23040 41530 23060 41690
rect 22980 41510 23060 41530
rect 23090 41690 23160 41710
rect 23090 41530 23110 41690
rect 23150 41530 23160 41690
rect 23090 41510 23160 41530
rect 23380 41550 23450 41570
rect 23380 41390 23390 41550
rect 23430 41390 23450 41550
rect 23380 41370 23450 41390
rect 23480 41550 23550 41570
rect 23480 41390 23500 41550
rect 23540 41390 23550 41550
rect 23480 41370 23550 41390
rect 5949 41160 6019 41180
rect 5949 41000 5959 41160
rect 5999 41000 6019 41160
rect 5949 40980 6019 41000
rect 6049 41160 6119 41180
rect 6049 41000 6069 41160
rect 6109 41000 6119 41160
rect 6049 40980 6119 41000
rect 6179 41160 6249 41180
rect 6179 41000 6189 41160
rect 6229 41000 6249 41160
rect 6179 40980 6249 41000
rect 6279 41160 6359 41180
rect 6279 41000 6299 41160
rect 6339 41000 6359 41160
rect 6279 40980 6359 41000
rect 6389 41160 6459 41180
rect 6389 41000 6409 41160
rect 6449 41000 6459 41160
rect 6389 40980 6459 41000
rect 6519 41160 6589 41180
rect 6519 41000 6529 41160
rect 6569 41000 6589 41160
rect 6519 40980 6589 41000
rect 6619 41160 6699 41180
rect 6619 41000 6639 41160
rect 6679 41000 6699 41160
rect 6619 40980 6699 41000
rect 6729 41160 6809 41180
rect 6729 41000 6749 41160
rect 6789 41000 6809 41160
rect 6729 40980 6809 41000
rect 6839 41160 6919 41180
rect 6839 41000 6859 41160
rect 6899 41000 6919 41160
rect 6839 40980 6919 41000
rect 6949 41160 7019 41180
rect 6949 41000 6969 41160
rect 7009 41000 7019 41160
rect 6949 40980 7019 41000
rect 7079 41160 7149 41180
rect 7079 41000 7089 41160
rect 7129 41000 7149 41160
rect 7079 40980 7149 41000
rect 7179 41160 7259 41180
rect 7179 41000 7199 41160
rect 7239 41000 7259 41160
rect 7179 40980 7259 41000
rect 7289 41160 7369 41180
rect 7289 41000 7309 41160
rect 7349 41000 7369 41160
rect 7289 40980 7369 41000
rect 7399 41160 7479 41180
rect 7399 41000 7419 41160
rect 7459 41000 7479 41160
rect 7399 40980 7479 41000
rect 7509 41160 7589 41180
rect 7509 41000 7529 41160
rect 7569 41000 7589 41160
rect 7509 40980 7589 41000
rect 7619 41160 7699 41180
rect 7619 41000 7639 41160
rect 7679 41000 7699 41160
rect 7619 40980 7699 41000
rect 7729 41160 7809 41180
rect 7729 41000 7749 41160
rect 7789 41000 7809 41160
rect 7729 40980 7809 41000
rect 7839 41160 7919 41180
rect 7839 41000 7859 41160
rect 7899 41000 7919 41160
rect 7839 40980 7919 41000
rect 7949 41160 8019 41180
rect 7949 41000 7969 41160
rect 8009 41000 8019 41160
rect 7949 40980 8019 41000
rect 8139 41160 8209 41180
rect 8139 41000 8149 41160
rect 8189 41000 8209 41160
rect 8139 40980 8209 41000
rect 8239 41160 8319 41180
rect 8239 41000 8259 41160
rect 8299 41000 8319 41160
rect 8239 40980 8319 41000
rect 8349 41160 8429 41180
rect 8349 41000 8369 41160
rect 8409 41000 8429 41160
rect 8349 40980 8429 41000
rect 8459 41160 8539 41180
rect 8459 41000 8479 41160
rect 8519 41000 8539 41160
rect 8459 40980 8539 41000
rect 8569 41160 8649 41180
rect 8569 41000 8589 41160
rect 8629 41000 8649 41160
rect 8569 40980 8649 41000
rect 8679 41160 8759 41180
rect 8679 41000 8699 41160
rect 8739 41000 8759 41160
rect 8679 40980 8759 41000
rect 8789 41160 8869 41180
rect 8789 41000 8809 41160
rect 8849 41000 8869 41160
rect 8789 40980 8869 41000
rect 8899 41160 8979 41180
rect 8899 41000 8919 41160
rect 8959 41000 8979 41160
rect 8899 40980 8979 41000
rect 9009 41160 9089 41180
rect 9009 41000 9029 41160
rect 9069 41000 9089 41160
rect 9009 40980 9089 41000
rect 9119 41160 9199 41180
rect 9119 41000 9139 41160
rect 9179 41000 9199 41160
rect 9119 40980 9199 41000
rect 9229 41160 9309 41180
rect 9229 41000 9249 41160
rect 9289 41000 9309 41160
rect 9229 40980 9309 41000
rect 9339 41160 9419 41180
rect 9339 41000 9359 41160
rect 9399 41000 9419 41160
rect 9339 40980 9419 41000
rect 9449 41160 9529 41180
rect 9449 41000 9469 41160
rect 9509 41000 9529 41160
rect 9449 40980 9529 41000
rect 9559 41160 9639 41180
rect 9559 41000 9579 41160
rect 9619 41000 9639 41160
rect 9559 40980 9639 41000
rect 9669 41160 9749 41180
rect 9669 41000 9689 41160
rect 9729 41000 9749 41160
rect 9669 40980 9749 41000
rect 9779 41160 9859 41180
rect 9779 41000 9799 41160
rect 9839 41000 9859 41160
rect 9779 40980 9859 41000
rect 9889 41160 9959 41180
rect 9889 41000 9909 41160
rect 9949 41000 9959 41160
rect 9889 40980 9959 41000
rect 2649 40540 2719 40560
rect 2649 39780 2659 40540
rect 2699 39780 2719 40540
rect 2649 39760 2719 39780
rect 2749 40540 2819 40560
rect 2749 39780 2769 40540
rect 2809 39780 2819 40540
rect 2749 39760 2819 39780
rect 2979 40540 3049 40560
rect 2979 39780 2989 40540
rect 3029 39780 3049 40540
rect 2979 39760 3049 39780
rect 3079 40540 3149 40560
rect 3079 39780 3099 40540
rect 3139 39780 3149 40540
rect 6349 39840 6419 39860
rect 3079 39760 3149 39780
rect 6349 39680 6359 39840
rect 6399 39680 6419 39840
rect 6349 39660 6419 39680
rect 6449 39840 6529 39860
rect 6449 39680 6469 39840
rect 6509 39680 6529 39840
rect 6449 39660 6529 39680
rect 6559 39840 6639 39860
rect 6559 39680 6579 39840
rect 6619 39680 6639 39840
rect 6559 39660 6639 39680
rect 6669 39840 6749 39860
rect 6669 39680 6689 39840
rect 6729 39680 6749 39840
rect 6669 39660 6749 39680
rect 6779 39840 6859 39860
rect 6779 39680 6799 39840
rect 6839 39680 6859 39840
rect 6779 39660 6859 39680
rect 6889 39840 6969 39860
rect 6889 39680 6909 39840
rect 6949 39680 6969 39840
rect 6889 39660 6969 39680
rect 6999 39840 7079 39860
rect 6999 39680 7019 39840
rect 7059 39680 7079 39840
rect 6999 39660 7079 39680
rect 7109 39840 7189 39860
rect 7109 39680 7129 39840
rect 7169 39680 7189 39840
rect 7109 39660 7189 39680
rect 7219 39840 7299 39860
rect 7219 39680 7239 39840
rect 7279 39680 7299 39840
rect 7219 39660 7299 39680
rect 7329 39840 7409 39860
rect 7329 39680 7349 39840
rect 7389 39680 7409 39840
rect 7329 39660 7409 39680
rect 7439 39840 7519 39860
rect 7439 39680 7459 39840
rect 7499 39680 7519 39840
rect 7439 39660 7519 39680
rect 7549 39840 7629 39860
rect 7549 39680 7569 39840
rect 7609 39680 7629 39840
rect 7549 39660 7629 39680
rect 7659 39840 7739 39860
rect 7659 39680 7679 39840
rect 7719 39680 7739 39840
rect 7659 39660 7739 39680
rect 7769 39840 7849 39860
rect 7769 39680 7789 39840
rect 7829 39680 7849 39840
rect 7769 39660 7849 39680
rect 7879 39840 7959 39860
rect 7879 39680 7899 39840
rect 7939 39680 7959 39840
rect 7879 39660 7959 39680
rect 7989 39840 8069 39860
rect 7989 39680 8009 39840
rect 8049 39680 8069 39840
rect 7989 39660 8069 39680
rect 8099 39840 8179 39860
rect 8099 39680 8119 39840
rect 8159 39680 8179 39840
rect 8099 39660 8179 39680
rect 8209 39840 8289 39860
rect 8209 39680 8229 39840
rect 8269 39680 8289 39840
rect 8209 39660 8289 39680
rect 8319 39840 8399 39860
rect 8319 39680 8339 39840
rect 8379 39680 8399 39840
rect 8319 39660 8399 39680
rect 8429 39840 8509 39860
rect 8429 39680 8449 39840
rect 8489 39680 8509 39840
rect 8429 39660 8509 39680
rect 8539 39840 8619 39860
rect 8539 39680 8559 39840
rect 8599 39680 8619 39840
rect 8539 39660 8619 39680
rect 8649 39840 8729 39860
rect 8649 39680 8669 39840
rect 8709 39680 8729 39840
rect 8649 39660 8729 39680
rect 8759 39840 8839 39860
rect 8759 39680 8779 39840
rect 8819 39680 8839 39840
rect 8759 39660 8839 39680
rect 8869 39840 8949 39860
rect 8869 39680 8889 39840
rect 8929 39680 8949 39840
rect 8869 39660 8949 39680
rect 8979 39840 9059 39860
rect 8979 39680 8999 39840
rect 9039 39680 9059 39840
rect 8979 39660 9059 39680
rect 9089 39840 9169 39860
rect 9089 39680 9109 39840
rect 9149 39680 9169 39840
rect 9089 39660 9169 39680
rect 9199 39840 9279 39860
rect 9199 39680 9219 39840
rect 9259 39680 9279 39840
rect 9199 39660 9279 39680
rect 9309 39840 9389 39860
rect 9309 39680 9329 39840
rect 9369 39680 9389 39840
rect 9309 39660 9389 39680
rect 9419 39840 9499 39860
rect 9419 39680 9439 39840
rect 9479 39680 9499 39840
rect 9419 39660 9499 39680
rect 9529 39840 9609 39860
rect 9529 39680 9549 39840
rect 9589 39680 9609 39840
rect 9529 39660 9609 39680
rect 9639 39840 9719 39860
rect 9639 39680 9659 39840
rect 9699 39680 9719 39840
rect 9639 39660 9719 39680
rect 9749 39840 9829 39860
rect 9749 39680 9769 39840
rect 9809 39680 9829 39840
rect 9749 39660 9829 39680
rect 9859 39840 9929 39860
rect 9859 39680 9879 39840
rect 9919 39680 9929 39840
rect 9859 39660 9929 39680
rect 3770 37030 3840 37050
rect 3770 36270 3780 37030
rect 3820 36270 3840 37030
rect 3770 36250 3840 36270
rect 3870 37030 3950 37050
rect 3870 36270 3890 37030
rect 3930 36270 3950 37030
rect 3870 36250 3950 36270
rect 3980 37030 4060 37050
rect 3980 36270 4000 37030
rect 4040 36270 4060 37030
rect 3980 36250 4060 36270
rect 4090 37030 4170 37050
rect 4090 36270 4110 37030
rect 4150 36270 4170 37030
rect 4090 36250 4170 36270
rect 4200 37030 4280 37050
rect 4200 36270 4220 37030
rect 4260 36270 4280 37030
rect 4200 36250 4280 36270
rect 4310 37030 4390 37050
rect 4310 36270 4330 37030
rect 4370 36270 4390 37030
rect 4310 36250 4390 36270
rect 4420 37030 4650 37050
rect 4420 36270 4510 37030
rect 4550 36270 4650 37030
rect 4420 36250 4650 36270
rect 4680 37030 4760 37050
rect 4680 36270 4700 37030
rect 4740 36270 4760 37030
rect 4680 36250 4760 36270
rect 4790 37030 4870 37050
rect 4790 36270 4810 37030
rect 4850 36270 4870 37030
rect 4790 36250 4870 36270
rect 4900 37030 4980 37050
rect 4900 36270 4920 37030
rect 4960 36270 4980 37030
rect 4900 36250 4980 36270
rect 5010 37030 5090 37050
rect 5010 36270 5030 37030
rect 5070 36270 5090 37030
rect 5010 36250 5090 36270
rect 5120 37030 5200 37050
rect 5120 36270 5140 37030
rect 5180 36270 5200 37030
rect 5120 36250 5200 36270
rect 5230 37030 5300 37050
rect 5230 36270 5250 37030
rect 5290 36270 5300 37030
rect 5460 37030 5530 37050
rect 5460 36670 5470 37030
rect 5510 36670 5530 37030
rect 5460 36650 5530 36670
rect 5560 37030 5640 37050
rect 5560 36670 5580 37030
rect 5620 36670 5640 37030
rect 5560 36650 5640 36670
rect 5670 37030 5750 37050
rect 5670 36670 5690 37030
rect 5730 36670 5750 37030
rect 5670 36650 5750 36670
rect 5780 37030 5860 37050
rect 5780 36670 5800 37030
rect 5840 36670 5860 37030
rect 5780 36650 5860 36670
rect 5890 37030 5970 37050
rect 5890 36670 5910 37030
rect 5950 36670 5970 37030
rect 5890 36650 5970 36670
rect 6000 37030 6080 37050
rect 6000 36670 6020 37030
rect 6060 36670 6080 37030
rect 6000 36650 6080 36670
rect 6110 37030 6180 37050
rect 6110 36670 6130 37030
rect 6170 36670 6180 37030
rect 6110 36650 6180 36670
rect 5230 36250 5300 36270
rect 6340 36570 6410 36590
rect 6340 36410 6350 36570
rect 6390 36410 6410 36570
rect 6340 36390 6410 36410
rect 6440 36570 6520 36590
rect 6440 36410 6460 36570
rect 6500 36410 6520 36570
rect 6440 36390 6520 36410
rect 6550 36570 6620 36590
rect 6550 36410 6570 36570
rect 6610 36410 6620 36570
rect 6550 36390 6620 36410
rect 6700 36190 6770 36590
rect 6800 36570 6880 36590
rect 6800 36210 6820 36570
rect 6860 36210 6880 36570
rect 6800 36190 6880 36210
rect 6910 36190 7030 36590
rect 7060 36570 7140 36590
rect 7060 36210 7080 36570
rect 7120 36210 7140 36570
rect 7060 36190 7140 36210
rect 7170 36190 7240 36590
rect 7300 36570 7370 36590
rect 7300 36410 7310 36570
rect 7350 36410 7370 36570
rect 7300 36390 7370 36410
rect 7400 36570 7480 36590
rect 7400 36410 7420 36570
rect 7460 36410 7480 36570
rect 7400 36390 7480 36410
rect 7510 36570 7580 36590
rect 7510 36410 7530 36570
rect 7570 36410 7580 36570
rect 7510 36390 7580 36410
rect 7680 36570 7750 36590
rect 7680 36410 7690 36570
rect 7730 36410 7750 36570
rect 7680 36390 7750 36410
rect 7780 36570 7860 36590
rect 7780 36410 7800 36570
rect 7840 36410 7860 36570
rect 7780 36390 7860 36410
rect 7890 36570 7960 36590
rect 7890 36410 7910 36570
rect 7950 36410 7960 36570
rect 7890 36390 7960 36410
rect 8060 36570 8130 36590
rect 8060 36410 8070 36570
rect 8110 36410 8130 36570
rect 8060 36390 8130 36410
rect 8160 36570 8240 36590
rect 8160 36410 8180 36570
rect 8220 36410 8240 36570
rect 8160 36390 8240 36410
rect 8270 36570 8340 36590
rect 8270 36410 8290 36570
rect 8330 36410 8340 36570
rect 8270 36390 8340 36410
rect 8440 36570 8510 36590
rect 8440 36410 8450 36570
rect 8490 36410 8510 36570
rect 8440 36390 8510 36410
rect 8540 36570 8620 36590
rect 8540 36410 8560 36570
rect 8600 36410 8620 36570
rect 8540 36390 8620 36410
rect 8650 36570 8720 36590
rect 8650 36410 8670 36570
rect 8710 36410 8720 36570
rect 8650 36390 8720 36410
rect 8780 36190 8850 36590
rect 8880 36570 8960 36590
rect 8880 36210 8900 36570
rect 8940 36210 8960 36570
rect 8880 36190 8960 36210
rect 8990 36190 9110 36590
rect 9140 36570 9220 36590
rect 9140 36210 9160 36570
rect 9200 36210 9220 36570
rect 9140 36190 9220 36210
rect 9250 36190 9320 36590
rect 9380 36570 9450 36590
rect 9380 36410 9390 36570
rect 9430 36410 9450 36570
rect 9380 36390 9450 36410
rect 9480 36570 9560 36590
rect 9480 36410 9500 36570
rect 9540 36410 9560 36570
rect 9480 36390 9560 36410
rect 9590 36570 9660 36590
rect 9590 36410 9610 36570
rect 9650 36410 9660 36570
rect 9590 36390 9660 36410
rect 9760 36570 9830 36590
rect 9760 36410 9770 36570
rect 9810 36410 9830 36570
rect 9760 36390 9830 36410
rect 9860 36570 9940 36590
rect 9860 36410 9880 36570
rect 9920 36410 9940 36570
rect 9860 36390 9940 36410
rect 9970 36570 10040 36590
rect 9970 36410 9990 36570
rect 10030 36410 10040 36570
rect 9970 36390 10040 36410
rect 10140 36570 10210 36590
rect 10140 36410 10150 36570
rect 10190 36410 10210 36570
rect 10140 36390 10210 36410
rect 10240 36570 10320 36590
rect 10240 36410 10260 36570
rect 10300 36410 10320 36570
rect 10240 36390 10320 36410
rect 10350 36570 10420 36590
rect 10350 36410 10370 36570
rect 10410 36410 10420 36570
rect 10350 36390 10420 36410
rect 10520 36570 10590 36590
rect 10520 36410 10530 36570
rect 10570 36410 10590 36570
rect 10520 36390 10590 36410
rect 10620 36570 10700 36590
rect 10620 36410 10640 36570
rect 10680 36410 10700 36570
rect 10620 36390 10700 36410
rect 10730 36570 10800 36590
rect 10730 36410 10750 36570
rect 10790 36410 10800 36570
rect 10730 36390 10800 36410
rect 16460 35820 16530 35840
rect 16460 35630 16470 35820
rect 16510 35630 16530 35820
rect 16460 35610 16530 35630
rect 16560 35820 16640 35840
rect 16560 35630 16580 35820
rect 16620 35630 16640 35820
rect 16560 35610 16640 35630
rect 16670 35820 16750 35840
rect 16670 35630 16690 35820
rect 16730 35630 16750 35820
rect 16670 35610 16750 35630
rect 16780 35820 16860 35840
rect 16780 35630 16800 35820
rect 16840 35630 16860 35820
rect 16780 35610 16860 35630
rect 16890 35820 16970 35840
rect 16890 35630 16910 35820
rect 16950 35630 16970 35820
rect 16890 35610 16970 35630
rect 17000 35820 17080 35840
rect 17000 35630 17020 35820
rect 17060 35630 17080 35820
rect 17000 35610 17080 35630
rect 17110 35820 17180 35840
rect 17110 35630 17130 35820
rect 17170 35630 17180 35820
rect 17110 35610 17180 35630
rect 16460 35330 16530 35350
rect 16460 34470 16470 35330
rect 16510 34470 16530 35330
rect 16460 34450 16530 34470
rect 16560 35330 16640 35350
rect 16560 34470 16580 35330
rect 16620 34470 16640 35330
rect 16560 34450 16640 34470
rect 16670 35330 16750 35350
rect 16670 34470 16690 35330
rect 16730 34470 16750 35330
rect 16670 34450 16750 34470
rect 16780 35330 16860 35350
rect 16780 34470 16800 35330
rect 16840 34470 16860 35330
rect 16780 34450 16860 34470
rect 16890 35330 16970 35350
rect 16890 34470 16910 35330
rect 16950 34470 16970 35330
rect 16890 34450 16970 34470
rect 17000 35330 17080 35350
rect 17000 34470 17020 35330
rect 17060 34470 17080 35330
rect 17000 34450 17080 34470
rect 17110 35330 17180 35350
rect 17110 34470 17130 35330
rect 17170 34470 17180 35330
rect 17350 35140 17420 35160
rect 17350 34980 17360 35140
rect 17400 34980 17420 35140
rect 17350 34960 17420 34980
rect 17450 35140 17520 35160
rect 17450 34980 17470 35140
rect 17510 34980 17520 35140
rect 18290 35140 18360 35160
rect 17450 34960 17520 34980
rect 17750 35090 17820 35110
rect 17750 34930 17760 35090
rect 17800 34930 17820 35090
rect 17750 34910 17820 34930
rect 17850 35090 17920 35110
rect 17850 34930 17870 35090
rect 17910 34930 17920 35090
rect 18290 34980 18300 35140
rect 18340 34980 18360 35140
rect 18290 34960 18360 34980
rect 18390 35140 18460 35160
rect 18390 34980 18410 35140
rect 18450 34980 18460 35140
rect 18390 34960 18460 34980
rect 18690 35140 18760 35160
rect 18690 34980 18700 35140
rect 18740 34980 18760 35140
rect 18690 34960 18760 34980
rect 18790 35140 18860 35160
rect 18790 34980 18810 35140
rect 18850 34980 18860 35140
rect 19760 35130 19830 35150
rect 18790 34960 18860 34980
rect 17850 34910 17920 34930
rect 19760 34970 19770 35130
rect 19810 34970 19830 35130
rect 19760 34950 19830 34970
rect 19860 35130 19930 35150
rect 19860 34970 19880 35130
rect 19920 34970 19930 35130
rect 19860 34950 19930 34970
rect 20010 35130 20080 35150
rect 20010 34970 20020 35130
rect 20060 34970 20080 35130
rect 20010 34950 20080 34970
rect 20110 35130 20180 35150
rect 20110 34970 20130 35130
rect 20170 34970 20180 35130
rect 21420 35820 21490 35840
rect 21420 35630 21430 35820
rect 21470 35630 21490 35820
rect 21420 35610 21490 35630
rect 21520 35820 21600 35840
rect 21520 35630 21540 35820
rect 21580 35630 21600 35820
rect 21520 35610 21600 35630
rect 21630 35820 21710 35840
rect 21630 35630 21650 35820
rect 21690 35630 21710 35820
rect 21630 35610 21710 35630
rect 21740 35820 21820 35840
rect 21740 35630 21760 35820
rect 21800 35630 21820 35820
rect 21740 35610 21820 35630
rect 21850 35820 21930 35840
rect 21850 35630 21870 35820
rect 21910 35630 21930 35820
rect 21850 35610 21930 35630
rect 21960 35820 22040 35840
rect 21960 35630 21980 35820
rect 22020 35630 22040 35820
rect 21960 35610 22040 35630
rect 22070 35820 22140 35840
rect 22070 35630 22090 35820
rect 22130 35630 22140 35820
rect 22070 35610 22140 35630
rect 21420 35330 21490 35350
rect 20110 34950 20180 34970
rect 19300 34830 19370 34850
rect 17110 34450 17180 34470
rect 17570 34620 17640 34640
rect 17570 34460 17580 34620
rect 17620 34460 17640 34620
rect 17570 34440 17640 34460
rect 17670 34620 17740 34640
rect 17670 34460 17690 34620
rect 17730 34460 17740 34620
rect 17670 34440 17740 34460
rect 18030 34620 18100 34640
rect 18030 34460 18040 34620
rect 18080 34460 18100 34620
rect 18030 34440 18100 34460
rect 18130 34620 18200 34640
rect 18130 34460 18150 34620
rect 18190 34460 18200 34620
rect 18130 34440 18200 34460
rect 18510 34620 18580 34640
rect 18510 34460 18520 34620
rect 18560 34460 18580 34620
rect 18510 34440 18580 34460
rect 18610 34620 18680 34640
rect 18610 34460 18630 34620
rect 18670 34460 18680 34620
rect 18610 34440 18680 34460
rect 18970 34620 19040 34640
rect 18970 34460 18980 34620
rect 19020 34460 19040 34620
rect 18970 34440 19040 34460
rect 19070 34620 19140 34640
rect 19070 34460 19090 34620
rect 19130 34460 19140 34620
rect 19070 34440 19140 34460
rect 19300 34470 19310 34830
rect 19350 34470 19370 34830
rect 19300 34450 19370 34470
rect 19400 34830 19470 34850
rect 19400 34470 19420 34830
rect 19460 34470 19470 34830
rect 21030 34830 21100 34850
rect 19400 34450 19470 34470
rect 19760 34550 19830 34570
rect 19760 34390 19770 34550
rect 19810 34390 19830 34550
rect 19760 34370 19830 34390
rect 19860 34550 19930 34570
rect 19860 34390 19880 34550
rect 19920 34390 19930 34550
rect 21030 34470 21040 34830
rect 21080 34470 21100 34830
rect 21030 34450 21100 34470
rect 21130 34830 21200 34850
rect 21130 34470 21150 34830
rect 21190 34470 21200 34830
rect 21130 34450 21200 34470
rect 21420 34470 21430 35330
rect 21470 34470 21490 35330
rect 21420 34450 21490 34470
rect 21520 35330 21600 35350
rect 21520 34470 21540 35330
rect 21580 34470 21600 35330
rect 21520 34450 21600 34470
rect 21630 35330 21710 35350
rect 21630 34470 21650 35330
rect 21690 34470 21710 35330
rect 21630 34450 21710 34470
rect 21740 35330 21820 35350
rect 21740 34470 21760 35330
rect 21800 34470 21820 35330
rect 21740 34450 21820 34470
rect 21850 35330 21930 35350
rect 21850 34470 21870 35330
rect 21910 34470 21930 35330
rect 21850 34450 21930 34470
rect 21960 35330 22040 35350
rect 21960 34470 21980 35330
rect 22020 34470 22040 35330
rect 21960 34450 22040 34470
rect 22070 35330 22140 35350
rect 22070 34470 22090 35330
rect 22130 34470 22140 35330
rect 22310 35140 22380 35160
rect 22310 34980 22320 35140
rect 22360 34980 22380 35140
rect 22310 34960 22380 34980
rect 22410 35140 22480 35160
rect 22410 34980 22430 35140
rect 22470 34980 22480 35140
rect 23250 35140 23320 35160
rect 22410 34960 22480 34980
rect 22710 35090 22780 35110
rect 22710 34930 22720 35090
rect 22760 34930 22780 35090
rect 22710 34910 22780 34930
rect 22810 35090 22880 35110
rect 22810 34930 22830 35090
rect 22870 34930 22880 35090
rect 23250 34980 23260 35140
rect 23300 34980 23320 35140
rect 23250 34960 23320 34980
rect 23350 35140 23420 35160
rect 23350 34980 23370 35140
rect 23410 34980 23420 35140
rect 23350 34960 23420 34980
rect 23650 35140 23720 35160
rect 23650 34980 23660 35140
rect 23700 34980 23720 35140
rect 23650 34960 23720 34980
rect 23750 35140 23820 35160
rect 23750 34980 23770 35140
rect 23810 34980 23820 35140
rect 24720 35130 24790 35150
rect 23750 34960 23820 34980
rect 22810 34910 22880 34930
rect 24720 34970 24730 35130
rect 24770 34970 24790 35130
rect 24720 34950 24790 34970
rect 24820 35130 24890 35150
rect 24820 34970 24840 35130
rect 24880 34970 24890 35130
rect 24820 34950 24890 34970
rect 24970 35130 25040 35150
rect 24970 34970 24980 35130
rect 25020 34970 25040 35130
rect 24970 34950 25040 34970
rect 25070 35130 25140 35150
rect 25070 34970 25090 35130
rect 25130 34970 25140 35130
rect 25070 34950 25140 34970
rect 24260 34830 24330 34850
rect 22070 34450 22140 34470
rect 22530 34620 22600 34640
rect 22530 34460 22540 34620
rect 22580 34460 22600 34620
rect 22530 34440 22600 34460
rect 22630 34620 22700 34640
rect 22630 34460 22650 34620
rect 22690 34460 22700 34620
rect 22630 34440 22700 34460
rect 22990 34620 23060 34640
rect 22990 34460 23000 34620
rect 23040 34460 23060 34620
rect 22990 34440 23060 34460
rect 23090 34620 23160 34640
rect 23090 34460 23110 34620
rect 23150 34460 23160 34620
rect 23090 34440 23160 34460
rect 23470 34620 23540 34640
rect 23470 34460 23480 34620
rect 23520 34460 23540 34620
rect 23470 34440 23540 34460
rect 23570 34620 23640 34640
rect 23570 34460 23590 34620
rect 23630 34460 23640 34620
rect 23570 34440 23640 34460
rect 23930 34620 24000 34640
rect 23930 34460 23940 34620
rect 23980 34460 24000 34620
rect 23930 34440 24000 34460
rect 24030 34620 24100 34640
rect 24030 34460 24050 34620
rect 24090 34460 24100 34620
rect 24030 34440 24100 34460
rect 24260 34470 24270 34830
rect 24310 34470 24330 34830
rect 24260 34450 24330 34470
rect 24360 34830 24430 34850
rect 24360 34470 24380 34830
rect 24420 34470 24430 34830
rect 24360 34450 24430 34470
rect 24720 34550 24790 34570
rect 19860 34370 19930 34390
rect 24720 34390 24730 34550
rect 24770 34390 24790 34550
rect 24720 34370 24790 34390
rect 24820 34550 24890 34570
rect 24820 34390 24840 34550
rect 24880 34390 24890 34550
rect 24820 34370 24890 34390
rect 16460 31760 16530 31780
rect 14108 31640 14178 31660
rect 2170 31580 2240 31600
rect 2170 30820 2180 31580
rect 2220 30820 2240 31580
rect 2170 30800 2240 30820
rect 2270 31580 2350 31600
rect 2270 30820 2290 31580
rect 2330 30820 2350 31580
rect 2270 30800 2350 30820
rect 2380 31580 2460 31600
rect 2380 30820 2400 31580
rect 2440 30820 2460 31580
rect 2380 30800 2460 30820
rect 2490 31580 2570 31600
rect 2490 30820 2510 31580
rect 2550 30820 2570 31580
rect 2490 30800 2570 30820
rect 2600 31580 2680 31600
rect 2600 30820 2620 31580
rect 2660 30820 2680 31580
rect 2600 30800 2680 30820
rect 2710 31580 2790 31600
rect 2710 30820 2730 31580
rect 2770 30820 2790 31580
rect 2710 30800 2790 30820
rect 2820 31580 3050 31600
rect 2820 30820 2910 31580
rect 2950 30820 3050 31580
rect 2820 30800 3050 30820
rect 3080 31580 3160 31600
rect 3080 30820 3100 31580
rect 3140 30820 3160 31580
rect 3080 30800 3160 30820
rect 3190 31580 3270 31600
rect 3190 30820 3210 31580
rect 3250 30820 3270 31580
rect 3190 30800 3270 30820
rect 3300 31580 3380 31600
rect 3300 30820 3320 31580
rect 3360 30820 3380 31580
rect 3300 30800 3380 30820
rect 3410 31580 3490 31600
rect 3410 30820 3430 31580
rect 3470 30820 3490 31580
rect 3410 30800 3490 30820
rect 3520 31580 3600 31600
rect 3520 30820 3540 31580
rect 3580 30820 3600 31580
rect 3520 30800 3600 30820
rect 3630 31580 3700 31600
rect 3630 30820 3650 31580
rect 3690 30820 3700 31580
rect 3860 31580 3930 31600
rect 3860 31220 3870 31580
rect 3910 31220 3930 31580
rect 3860 31200 3930 31220
rect 3960 31580 4040 31600
rect 3960 31220 3980 31580
rect 4020 31220 4040 31580
rect 3960 31200 4040 31220
rect 4070 31580 4150 31600
rect 4070 31220 4090 31580
rect 4130 31220 4150 31580
rect 4070 31200 4150 31220
rect 4180 31580 4260 31600
rect 4180 31220 4200 31580
rect 4240 31220 4260 31580
rect 4180 31200 4260 31220
rect 4290 31580 4370 31600
rect 4290 31220 4310 31580
rect 4350 31220 4370 31580
rect 4290 31200 4370 31220
rect 4400 31580 4480 31600
rect 4400 31220 4420 31580
rect 4460 31220 4480 31580
rect 4400 31200 4480 31220
rect 4510 31580 4580 31600
rect 4510 31220 4530 31580
rect 4570 31220 4580 31580
rect 4510 31200 4580 31220
rect 4720 31580 4790 31600
rect 4720 31220 4730 31580
rect 4770 31220 4790 31580
rect 4720 31200 4790 31220
rect 4820 31580 4900 31600
rect 4820 31220 4840 31580
rect 4880 31220 4900 31580
rect 4820 31200 4900 31220
rect 4930 31580 5010 31600
rect 4930 31220 4950 31580
rect 4990 31220 5010 31580
rect 4930 31200 5010 31220
rect 5040 31580 5120 31600
rect 5040 31220 5060 31580
rect 5100 31220 5120 31580
rect 5040 31200 5120 31220
rect 5150 31580 5230 31600
rect 5150 31220 5170 31580
rect 5210 31220 5230 31580
rect 5150 31200 5230 31220
rect 5260 31580 5340 31600
rect 5260 31220 5280 31580
rect 5320 31220 5340 31580
rect 5260 31200 5340 31220
rect 5370 31580 5440 31600
rect 5370 31220 5390 31580
rect 5430 31220 5440 31580
rect 5370 31200 5440 31220
rect 5580 31580 5650 31600
rect 5580 31220 5590 31580
rect 5630 31220 5650 31580
rect 5580 31200 5650 31220
rect 5680 31580 5760 31600
rect 5680 31220 5700 31580
rect 5740 31220 5760 31580
rect 5680 31200 5760 31220
rect 5790 31580 5870 31600
rect 5790 31220 5810 31580
rect 5850 31220 5870 31580
rect 5790 31200 5870 31220
rect 5900 31580 5980 31600
rect 5900 31220 5920 31580
rect 5960 31220 5980 31580
rect 5900 31200 5980 31220
rect 6010 31580 6090 31600
rect 6010 31220 6030 31580
rect 6070 31220 6090 31580
rect 6010 31200 6090 31220
rect 6120 31580 6200 31600
rect 6120 31220 6140 31580
rect 6180 31220 6200 31580
rect 6120 31200 6200 31220
rect 6230 31580 6300 31600
rect 6230 31220 6250 31580
rect 6290 31220 6300 31580
rect 14108 31380 14118 31640
rect 14158 31380 14178 31640
rect 14108 31360 14178 31380
rect 14208 31640 14278 31660
rect 14208 31380 14228 31640
rect 14268 31380 14278 31640
rect 16460 31570 16470 31760
rect 16510 31570 16530 31760
rect 16460 31550 16530 31570
rect 16560 31760 16640 31780
rect 16560 31570 16580 31760
rect 16620 31570 16640 31760
rect 16560 31550 16640 31570
rect 16670 31760 16750 31780
rect 16670 31570 16690 31760
rect 16730 31570 16750 31760
rect 16670 31550 16750 31570
rect 16780 31760 16860 31780
rect 16780 31570 16800 31760
rect 16840 31570 16860 31760
rect 16780 31550 16860 31570
rect 16890 31760 16970 31780
rect 16890 31570 16910 31760
rect 16950 31570 16970 31760
rect 16890 31550 16970 31570
rect 17000 31760 17080 31780
rect 17000 31570 17020 31760
rect 17060 31570 17080 31760
rect 17000 31550 17080 31570
rect 17110 31760 17180 31780
rect 17110 31570 17130 31760
rect 17170 31570 17180 31760
rect 17110 31550 17180 31570
rect 14208 31360 14278 31380
rect 16460 31270 16530 31290
rect 6230 31200 6300 31220
rect 6400 31220 6470 31240
rect 3630 30800 3700 30820
rect 6400 31060 6410 31220
rect 6450 31060 6470 31220
rect 6400 31040 6470 31060
rect 6500 31220 6580 31240
rect 6500 31060 6520 31220
rect 6560 31060 6580 31220
rect 6500 31040 6580 31060
rect 6610 31220 6680 31240
rect 6610 31060 6630 31220
rect 6670 31060 6680 31220
rect 6610 31040 6680 31060
rect 6760 30840 6830 31240
rect 6860 31220 6940 31240
rect 6860 30860 6880 31220
rect 6920 30860 6940 31220
rect 6860 30840 6940 30860
rect 6970 30840 7090 31240
rect 7120 31220 7200 31240
rect 7120 30860 7140 31220
rect 7180 30860 7200 31220
rect 7120 30840 7200 30860
rect 7230 30840 7300 31240
rect 7360 31220 7430 31240
rect 7360 31060 7370 31220
rect 7410 31060 7430 31220
rect 7360 31040 7430 31060
rect 7460 31220 7540 31240
rect 7460 31060 7480 31220
rect 7520 31060 7540 31220
rect 7460 31040 7540 31060
rect 7570 31220 7640 31240
rect 7570 31060 7590 31220
rect 7630 31060 7640 31220
rect 7570 31040 7640 31060
rect 7740 31220 7810 31240
rect 7740 31060 7750 31220
rect 7790 31060 7810 31220
rect 7740 31040 7810 31060
rect 7840 31220 7920 31240
rect 7840 31060 7860 31220
rect 7900 31060 7920 31220
rect 7840 31040 7920 31060
rect 7950 31220 8020 31240
rect 7950 31060 7970 31220
rect 8010 31060 8020 31220
rect 7950 31040 8020 31060
rect 8120 31220 8190 31240
rect 8120 31060 8130 31220
rect 8170 31060 8190 31220
rect 8120 31040 8190 31060
rect 8220 31220 8300 31240
rect 8220 31060 8240 31220
rect 8280 31060 8300 31220
rect 8220 31040 8300 31060
rect 8330 31220 8400 31240
rect 8330 31060 8350 31220
rect 8390 31060 8400 31220
rect 8330 31040 8400 31060
rect 8500 31220 8570 31240
rect 8500 31060 8510 31220
rect 8550 31060 8570 31220
rect 8500 31040 8570 31060
rect 8600 31220 8680 31240
rect 8600 31060 8620 31220
rect 8660 31060 8680 31220
rect 8600 31040 8680 31060
rect 8710 31220 8780 31240
rect 8710 31060 8730 31220
rect 8770 31060 8780 31220
rect 8710 31040 8780 31060
rect 8840 30840 8910 31240
rect 8940 31220 9020 31240
rect 8940 30860 8960 31220
rect 9000 30860 9020 31220
rect 8940 30840 9020 30860
rect 9050 30840 9170 31240
rect 9200 31220 9280 31240
rect 9200 30860 9220 31220
rect 9260 30860 9280 31220
rect 9200 30840 9280 30860
rect 9310 30840 9380 31240
rect 9440 31220 9510 31240
rect 9440 31060 9450 31220
rect 9490 31060 9510 31220
rect 9440 31040 9510 31060
rect 9540 31220 9620 31240
rect 9540 31060 9560 31220
rect 9600 31060 9620 31220
rect 9540 31040 9620 31060
rect 9650 31220 9720 31240
rect 9650 31060 9670 31220
rect 9710 31060 9720 31220
rect 9650 31040 9720 31060
rect 9820 31220 9890 31240
rect 9820 31060 9830 31220
rect 9870 31060 9890 31220
rect 9820 31040 9890 31060
rect 9920 31220 10000 31240
rect 9920 31060 9940 31220
rect 9980 31060 10000 31220
rect 9920 31040 10000 31060
rect 10030 31220 10100 31240
rect 10030 31060 10050 31220
rect 10090 31060 10100 31220
rect 10030 31040 10100 31060
rect 10200 31220 10270 31240
rect 10200 31060 10210 31220
rect 10250 31060 10270 31220
rect 10200 31040 10270 31060
rect 10300 31220 10380 31240
rect 10300 31060 10320 31220
rect 10360 31060 10380 31220
rect 10300 31040 10380 31060
rect 10410 31220 10480 31240
rect 10410 31060 10430 31220
rect 10470 31060 10480 31220
rect 10410 31040 10480 31060
rect 10580 31220 10650 31240
rect 10580 31060 10590 31220
rect 10630 31060 10650 31220
rect 10580 31040 10650 31060
rect 10680 31220 10760 31240
rect 10680 31060 10700 31220
rect 10740 31060 10760 31220
rect 10680 31040 10760 31060
rect 10790 31220 10860 31240
rect 10790 31060 10810 31220
rect 10850 31060 10860 31220
rect 10790 31040 10860 31060
rect 10960 31220 11030 31240
rect 10960 31060 10970 31220
rect 11010 31060 11030 31220
rect 10960 31040 11030 31060
rect 11060 31220 11140 31240
rect 11060 31060 11080 31220
rect 11120 31060 11140 31220
rect 11060 31040 11140 31060
rect 11170 31220 11240 31240
rect 11170 31060 11190 31220
rect 11230 31060 11240 31220
rect 11170 31040 11240 31060
rect 16460 30410 16470 31270
rect 16510 30410 16530 31270
rect 16460 30390 16530 30410
rect 16560 31270 16640 31290
rect 16560 30410 16580 31270
rect 16620 30410 16640 31270
rect 16560 30390 16640 30410
rect 16670 31270 16750 31290
rect 16670 30410 16690 31270
rect 16730 30410 16750 31270
rect 16670 30390 16750 30410
rect 16780 31270 16860 31290
rect 16780 30410 16800 31270
rect 16840 30410 16860 31270
rect 16780 30390 16860 30410
rect 16890 31270 16970 31290
rect 16890 30410 16910 31270
rect 16950 30410 16970 31270
rect 16890 30390 16970 30410
rect 17000 31270 17080 31290
rect 17000 30410 17020 31270
rect 17060 30410 17080 31270
rect 17000 30390 17080 30410
rect 17110 31270 17180 31290
rect 17110 30410 17130 31270
rect 17170 30410 17180 31270
rect 17350 31080 17420 31100
rect 17350 30920 17360 31080
rect 17400 30920 17420 31080
rect 17350 30900 17420 30920
rect 17450 31080 17520 31100
rect 17450 30920 17470 31080
rect 17510 30920 17520 31080
rect 18290 31080 18360 31100
rect 17450 30900 17520 30920
rect 17750 31030 17820 31050
rect 17750 30870 17760 31030
rect 17800 30870 17820 31030
rect 17750 30850 17820 30870
rect 17850 31030 17920 31050
rect 17850 30870 17870 31030
rect 17910 30870 17920 31030
rect 18290 30920 18300 31080
rect 18340 30920 18360 31080
rect 18290 30900 18360 30920
rect 18390 31080 18460 31100
rect 18390 30920 18410 31080
rect 18450 30920 18460 31080
rect 18390 30900 18460 30920
rect 18690 31080 18760 31100
rect 18690 30920 18700 31080
rect 18740 30920 18760 31080
rect 18690 30900 18760 30920
rect 18790 31080 18860 31100
rect 18790 30920 18810 31080
rect 18850 30920 18860 31080
rect 20020 31070 20090 31090
rect 18790 30900 18860 30920
rect 17850 30850 17920 30870
rect 20020 30910 20030 31070
rect 20070 30910 20090 31070
rect 20020 30890 20090 30910
rect 20120 31070 20190 31090
rect 20120 30910 20140 31070
rect 20180 30910 20190 31070
rect 20120 30890 20190 30910
rect 20270 31070 20340 31090
rect 20270 30910 20280 31070
rect 20320 30910 20340 31070
rect 20270 30890 20340 30910
rect 20370 31070 20440 31090
rect 20370 30910 20390 31070
rect 20430 30910 20440 31070
rect 21480 31750 21550 31770
rect 21480 31560 21490 31750
rect 21530 31560 21550 31750
rect 21480 31540 21550 31560
rect 21580 31750 21660 31770
rect 21580 31560 21600 31750
rect 21640 31560 21660 31750
rect 21580 31540 21660 31560
rect 21690 31750 21770 31770
rect 21690 31560 21710 31750
rect 21750 31560 21770 31750
rect 21690 31540 21770 31560
rect 21800 31750 21880 31770
rect 21800 31560 21820 31750
rect 21860 31560 21880 31750
rect 21800 31540 21880 31560
rect 21910 31750 21990 31770
rect 21910 31560 21930 31750
rect 21970 31560 21990 31750
rect 21910 31540 21990 31560
rect 22020 31750 22100 31770
rect 22020 31560 22040 31750
rect 22080 31560 22100 31750
rect 22020 31540 22100 31560
rect 22130 31750 22200 31770
rect 22130 31560 22150 31750
rect 22190 31560 22200 31750
rect 22130 31540 22200 31560
rect 21480 31260 21550 31280
rect 20370 30890 20440 30910
rect 19300 30770 19370 30790
rect 17110 30390 17180 30410
rect 17570 30560 17640 30580
rect 17570 30400 17580 30560
rect 17620 30400 17640 30560
rect 17570 30380 17640 30400
rect 17670 30560 17740 30580
rect 17670 30400 17690 30560
rect 17730 30400 17740 30560
rect 17670 30380 17740 30400
rect 18030 30560 18100 30580
rect 18030 30400 18040 30560
rect 18080 30400 18100 30560
rect 18030 30380 18100 30400
rect 18130 30560 18200 30580
rect 18130 30400 18150 30560
rect 18190 30400 18200 30560
rect 18130 30380 18200 30400
rect 18510 30560 18580 30580
rect 18510 30400 18520 30560
rect 18560 30400 18580 30560
rect 18510 30380 18580 30400
rect 18610 30560 18680 30580
rect 18610 30400 18630 30560
rect 18670 30400 18680 30560
rect 18610 30380 18680 30400
rect 18970 30560 19040 30580
rect 18970 30400 18980 30560
rect 19020 30400 19040 30560
rect 18970 30380 19040 30400
rect 19070 30560 19140 30580
rect 19070 30400 19090 30560
rect 19130 30400 19140 30560
rect 19070 30380 19140 30400
rect 19300 30410 19310 30770
rect 19350 30410 19370 30770
rect 19300 30390 19370 30410
rect 19400 30770 19470 30790
rect 19400 30410 19420 30770
rect 19460 30410 19470 30770
rect 19400 30390 19470 30410
rect 19560 30770 19630 30790
rect 19560 30410 19570 30770
rect 19610 30410 19630 30770
rect 19560 30390 19630 30410
rect 19660 30770 19730 30790
rect 19660 30410 19680 30770
rect 19720 30410 19730 30770
rect 21090 30770 21160 30790
rect 19660 30390 19730 30410
rect 20020 30490 20090 30510
rect 20020 30330 20030 30490
rect 20070 30330 20090 30490
rect 20020 30310 20090 30330
rect 20120 30490 20190 30510
rect 20120 30330 20140 30490
rect 20180 30330 20190 30490
rect 21090 30410 21100 30770
rect 21140 30410 21160 30770
rect 21090 30390 21160 30410
rect 21190 30770 21260 30790
rect 21190 30410 21210 30770
rect 21250 30410 21260 30770
rect 21190 30390 21260 30410
rect 21480 30400 21490 31260
rect 21530 30400 21550 31260
rect 21480 30380 21550 30400
rect 21580 31260 21660 31280
rect 21580 30400 21600 31260
rect 21640 30400 21660 31260
rect 21580 30380 21660 30400
rect 21690 31260 21770 31280
rect 21690 30400 21710 31260
rect 21750 30400 21770 31260
rect 21690 30380 21770 30400
rect 21800 31260 21880 31280
rect 21800 30400 21820 31260
rect 21860 30400 21880 31260
rect 21800 30380 21880 30400
rect 21910 31260 21990 31280
rect 21910 30400 21930 31260
rect 21970 30400 21990 31260
rect 21910 30380 21990 30400
rect 22020 31260 22100 31280
rect 22020 30400 22040 31260
rect 22080 30400 22100 31260
rect 22020 30380 22100 30400
rect 22130 31260 22200 31280
rect 22130 30400 22150 31260
rect 22190 30400 22200 31260
rect 22370 31070 22440 31090
rect 22370 30910 22380 31070
rect 22420 30910 22440 31070
rect 22370 30890 22440 30910
rect 22470 31070 22540 31090
rect 22470 30910 22490 31070
rect 22530 30910 22540 31070
rect 23310 31070 23380 31090
rect 22470 30890 22540 30910
rect 22770 31020 22840 31040
rect 22770 30860 22780 31020
rect 22820 30860 22840 31020
rect 22770 30840 22840 30860
rect 22870 31020 22940 31040
rect 22870 30860 22890 31020
rect 22930 30860 22940 31020
rect 23310 30910 23320 31070
rect 23360 30910 23380 31070
rect 23310 30890 23380 30910
rect 23410 31070 23480 31090
rect 23410 30910 23430 31070
rect 23470 30910 23480 31070
rect 23410 30890 23480 30910
rect 23710 31070 23780 31090
rect 23710 30910 23720 31070
rect 23760 30910 23780 31070
rect 23710 30890 23780 30910
rect 23810 31070 23880 31090
rect 23810 30910 23830 31070
rect 23870 30910 23880 31070
rect 24980 31060 25050 31080
rect 23810 30890 23880 30910
rect 22870 30840 22940 30860
rect 24980 30900 24990 31060
rect 25030 30900 25050 31060
rect 24980 30880 25050 30900
rect 25080 31060 25150 31080
rect 25080 30900 25100 31060
rect 25140 30900 25150 31060
rect 25080 30880 25150 30900
rect 25230 31060 25300 31080
rect 25230 30900 25240 31060
rect 25280 30900 25300 31060
rect 25230 30880 25300 30900
rect 25330 31060 25400 31080
rect 25330 30900 25350 31060
rect 25390 30900 25400 31060
rect 25330 30880 25400 30900
rect 24320 30760 24390 30780
rect 22130 30380 22200 30400
rect 22590 30550 22660 30570
rect 22590 30390 22600 30550
rect 22640 30390 22660 30550
rect 22590 30370 22660 30390
rect 22690 30550 22760 30570
rect 22690 30390 22710 30550
rect 22750 30390 22760 30550
rect 22690 30370 22760 30390
rect 23050 30550 23120 30570
rect 23050 30390 23060 30550
rect 23100 30390 23120 30550
rect 23050 30370 23120 30390
rect 23150 30550 23220 30570
rect 23150 30390 23170 30550
rect 23210 30390 23220 30550
rect 23150 30370 23220 30390
rect 23530 30550 23600 30570
rect 23530 30390 23540 30550
rect 23580 30390 23600 30550
rect 23530 30370 23600 30390
rect 23630 30550 23700 30570
rect 23630 30390 23650 30550
rect 23690 30390 23700 30550
rect 23630 30370 23700 30390
rect 23990 30550 24060 30570
rect 23990 30390 24000 30550
rect 24040 30390 24060 30550
rect 23990 30370 24060 30390
rect 24090 30550 24160 30570
rect 24090 30390 24110 30550
rect 24150 30390 24160 30550
rect 24090 30370 24160 30390
rect 24320 30400 24330 30760
rect 24370 30400 24390 30760
rect 24320 30380 24390 30400
rect 24420 30760 24490 30780
rect 24420 30400 24440 30760
rect 24480 30400 24490 30760
rect 24420 30380 24490 30400
rect 24580 30760 24650 30780
rect 24580 30400 24590 30760
rect 24630 30400 24650 30760
rect 24580 30380 24650 30400
rect 24680 30760 24750 30780
rect 24680 30400 24700 30760
rect 24740 30400 24750 30760
rect 24680 30380 24750 30400
rect 24980 30480 25050 30500
rect 20120 30310 20190 30330
rect 24980 30320 24990 30480
rect 25030 30320 25050 30480
rect 24980 30300 25050 30320
rect 25080 30480 25150 30500
rect 25080 30320 25100 30480
rect 25140 30320 25150 30480
rect 25080 30300 25150 30320
rect 8860 24810 8930 24830
rect 8480 24740 8550 24760
rect 7320 24550 7390 24570
rect 7320 24390 7330 24550
rect 7370 24390 7390 24550
rect 7320 24370 7390 24390
rect 7420 24550 7500 24570
rect 7420 24390 7440 24550
rect 7480 24390 7500 24550
rect 7420 24370 7500 24390
rect 7530 24550 7600 24570
rect 7530 24390 7550 24550
rect 7590 24390 7600 24550
rect 7530 24370 7600 24390
rect 7850 24550 7920 24570
rect 7850 24390 7860 24550
rect 7900 24390 7920 24550
rect 7850 24370 7920 24390
rect 7950 24550 8030 24570
rect 7950 24390 7970 24550
rect 8010 24390 8030 24550
rect 7950 24370 8030 24390
rect 8060 24550 8130 24570
rect 8060 24390 8080 24550
rect 8120 24390 8130 24550
rect 8060 24370 8130 24390
rect 8480 24380 8490 24740
rect 8530 24380 8550 24740
rect 8480 24360 8550 24380
rect 8580 24740 8700 24760
rect 8580 24380 8620 24740
rect 8660 24380 8700 24740
rect 8580 24360 8700 24380
rect 8730 24740 8800 24760
rect 8730 24380 8750 24740
rect 8790 24380 8800 24740
rect 8860 24650 8870 24810
rect 8910 24650 8930 24810
rect 8860 24630 8930 24650
rect 8960 24810 9030 24830
rect 8960 24650 8980 24810
rect 9020 24650 9030 24810
rect 8960 24630 9030 24650
rect 8730 24360 8800 24380
rect 9220 24540 9290 24560
rect 9220 24380 9230 24540
rect 9270 24380 9290 24540
rect 9220 24360 9290 24380
rect 9320 24540 9400 24560
rect 9320 24380 9340 24540
rect 9380 24380 9400 24540
rect 9320 24360 9400 24380
rect 9430 24540 9500 24560
rect 9430 24380 9450 24540
rect 9490 24380 9500 24540
rect 9430 24360 9500 24380
rect 9560 24360 9630 24760
rect 9660 24740 9740 24760
rect 9660 24380 9680 24740
rect 9720 24380 9740 24740
rect 9660 24360 9740 24380
rect 9770 24360 9890 24760
rect 9920 24740 10000 24760
rect 9920 24380 9940 24740
rect 9980 24380 10000 24740
rect 9920 24360 10000 24380
rect 10030 24360 10100 24760
rect 10160 24540 10230 24560
rect 10160 24380 10170 24540
rect 10210 24380 10230 24540
rect 10160 24360 10230 24380
rect 10260 24540 10340 24560
rect 10260 24380 10280 24540
rect 10320 24380 10340 24540
rect 10260 24360 10340 24380
rect 10370 24540 10440 24560
rect 10370 24380 10390 24540
rect 10430 24380 10440 24540
rect 10370 24360 10440 24380
rect 10550 24360 10620 24760
rect 10650 24740 10730 24760
rect 10650 24380 10670 24740
rect 10710 24380 10730 24740
rect 10650 24360 10730 24380
rect 10760 24360 10880 24760
rect 10910 24740 10990 24760
rect 10910 24380 10930 24740
rect 10970 24380 10990 24740
rect 10910 24360 10990 24380
rect 11020 24360 11090 24760
rect 11150 24540 11220 24560
rect 11150 24380 11160 24540
rect 11200 24380 11220 24540
rect 11150 24360 11220 24380
rect 11250 24540 11330 24560
rect 11250 24380 11270 24540
rect 11310 24380 11330 24540
rect 11250 24360 11330 24380
rect 11360 24540 11430 24560
rect 11360 24380 11380 24540
rect 11420 24380 11430 24540
rect 11360 24360 11430 24380
rect 11550 24360 11620 24760
rect 11650 24740 11730 24760
rect 11650 24380 11670 24740
rect 11710 24380 11730 24740
rect 11650 24360 11730 24380
rect 11760 24360 11880 24760
rect 11910 24740 11990 24760
rect 11910 24380 11930 24740
rect 11970 24380 11990 24740
rect 11910 24360 11990 24380
rect 12020 24360 12090 24760
rect 12880 24820 12950 24840
rect 12880 24660 12890 24820
rect 12930 24660 12950 24820
rect 12880 24640 12950 24660
rect 12980 24820 13050 24840
rect 12980 24660 13000 24820
rect 13040 24660 13050 24820
rect 12980 24640 13050 24660
rect 13110 24820 13180 24840
rect 13110 24660 13120 24820
rect 13160 24660 13180 24820
rect 13110 24640 13180 24660
rect 13210 24820 13290 24840
rect 13210 24660 13230 24820
rect 13270 24660 13290 24820
rect 13210 24640 13290 24660
rect 13320 24820 13390 24840
rect 13320 24660 13340 24820
rect 13380 24660 13390 24820
rect 13320 24640 13390 24660
rect 13450 24820 13520 24840
rect 13450 24660 13460 24820
rect 13500 24660 13520 24820
rect 13450 24640 13520 24660
rect 13550 24820 13630 24840
rect 13550 24660 13570 24820
rect 13610 24660 13630 24820
rect 13550 24640 13630 24660
rect 13660 24820 13740 24840
rect 13660 24660 13680 24820
rect 13720 24660 13740 24820
rect 13660 24640 13740 24660
rect 13770 24820 13850 24840
rect 13770 24660 13790 24820
rect 13830 24660 13850 24820
rect 13770 24640 13850 24660
rect 13880 24820 13950 24840
rect 13880 24660 13900 24820
rect 13940 24660 13950 24820
rect 13880 24640 13950 24660
rect 14010 24820 14080 24840
rect 14010 24660 14020 24820
rect 14060 24660 14080 24820
rect 14010 24640 14080 24660
rect 14110 24820 14190 24840
rect 14110 24660 14130 24820
rect 14170 24660 14190 24820
rect 14110 24640 14190 24660
rect 14220 24820 14300 24840
rect 14220 24660 14240 24820
rect 14280 24660 14300 24820
rect 14220 24640 14300 24660
rect 14330 24820 14410 24840
rect 14330 24660 14350 24820
rect 14390 24660 14410 24820
rect 14330 24640 14410 24660
rect 14440 24820 14520 24840
rect 14440 24660 14460 24820
rect 14500 24660 14520 24820
rect 14440 24640 14520 24660
rect 14550 24820 14630 24840
rect 14550 24660 14570 24820
rect 14610 24660 14630 24820
rect 14550 24640 14630 24660
rect 14660 24820 14740 24840
rect 14660 24660 14680 24820
rect 14720 24660 14740 24820
rect 14660 24640 14740 24660
rect 14770 24820 14850 24840
rect 14770 24660 14790 24820
rect 14830 24660 14850 24820
rect 14770 24640 14850 24660
rect 14880 24820 14950 24840
rect 14880 24660 14900 24820
rect 14940 24660 14950 24820
rect 14880 24640 14950 24660
rect 15070 24820 15140 24840
rect 15070 24660 15080 24820
rect 15120 24660 15140 24820
rect 15070 24640 15140 24660
rect 15170 24820 15250 24840
rect 15170 24660 15190 24820
rect 15230 24660 15250 24820
rect 15170 24640 15250 24660
rect 15280 24820 15360 24840
rect 15280 24660 15300 24820
rect 15340 24660 15360 24820
rect 15280 24640 15360 24660
rect 15390 24820 15470 24840
rect 15390 24660 15410 24820
rect 15450 24660 15470 24820
rect 15390 24640 15470 24660
rect 15500 24820 15580 24840
rect 15500 24660 15520 24820
rect 15560 24660 15580 24820
rect 15500 24640 15580 24660
rect 15610 24820 15690 24840
rect 15610 24660 15630 24820
rect 15670 24660 15690 24820
rect 15610 24640 15690 24660
rect 15720 24820 15800 24840
rect 15720 24660 15740 24820
rect 15780 24660 15800 24820
rect 15720 24640 15800 24660
rect 15830 24820 15910 24840
rect 15830 24660 15850 24820
rect 15890 24660 15910 24820
rect 15830 24640 15910 24660
rect 15940 24820 16020 24840
rect 15940 24660 15960 24820
rect 16000 24660 16020 24820
rect 15940 24640 16020 24660
rect 16050 24820 16130 24840
rect 16050 24660 16070 24820
rect 16110 24660 16130 24820
rect 16050 24640 16130 24660
rect 16160 24820 16240 24840
rect 16160 24660 16180 24820
rect 16220 24660 16240 24820
rect 16160 24640 16240 24660
rect 16270 24820 16350 24840
rect 16270 24660 16290 24820
rect 16330 24660 16350 24820
rect 16270 24640 16350 24660
rect 16380 24820 16460 24840
rect 16380 24660 16400 24820
rect 16440 24660 16460 24820
rect 16380 24640 16460 24660
rect 16490 24820 16570 24840
rect 16490 24660 16510 24820
rect 16550 24660 16570 24820
rect 16490 24640 16570 24660
rect 16600 24820 16680 24840
rect 16600 24660 16620 24820
rect 16660 24660 16680 24820
rect 16600 24640 16680 24660
rect 16710 24820 16790 24840
rect 16710 24660 16730 24820
rect 16770 24660 16790 24820
rect 16710 24640 16790 24660
rect 16820 24820 16890 24840
rect 16820 24660 16840 24820
rect 16880 24660 16890 24820
rect 16820 24640 16890 24660
rect 17020 24820 17090 24840
rect 17020 24660 17030 24820
rect 17070 24660 17090 24820
rect 17020 24640 17090 24660
rect 17120 24820 17200 24840
rect 17120 24660 17140 24820
rect 17180 24660 17200 24820
rect 17120 24640 17200 24660
rect 17230 24820 17310 24840
rect 17230 24660 17250 24820
rect 17290 24660 17310 24820
rect 17230 24640 17310 24660
rect 17340 24820 17420 24840
rect 17340 24660 17360 24820
rect 17400 24660 17420 24820
rect 17340 24640 17420 24660
rect 17450 24820 17530 24840
rect 17450 24660 17470 24820
rect 17510 24660 17530 24820
rect 17450 24640 17530 24660
rect 17560 24820 17640 24840
rect 17560 24660 17580 24820
rect 17620 24660 17640 24820
rect 17560 24640 17640 24660
rect 17670 24820 17750 24840
rect 17670 24660 17690 24820
rect 17730 24660 17750 24820
rect 17670 24640 17750 24660
rect 17780 24820 17860 24840
rect 17780 24660 17800 24820
rect 17840 24660 17860 24820
rect 17780 24640 17860 24660
rect 17890 24820 17970 24840
rect 17890 24660 17910 24820
rect 17950 24660 17970 24820
rect 17890 24640 17970 24660
rect 18000 24820 18080 24840
rect 18000 24660 18020 24820
rect 18060 24660 18080 24820
rect 18000 24640 18080 24660
rect 18110 24820 18190 24840
rect 18110 24660 18130 24820
rect 18170 24660 18190 24820
rect 18110 24640 18190 24660
rect 18220 24820 18300 24840
rect 18220 24660 18240 24820
rect 18280 24660 18300 24820
rect 18220 24640 18300 24660
rect 18330 24820 18410 24840
rect 18330 24660 18350 24820
rect 18390 24660 18410 24820
rect 18330 24640 18410 24660
rect 18440 24820 18520 24840
rect 18440 24660 18460 24820
rect 18500 24660 18520 24820
rect 18440 24640 18520 24660
rect 18550 24820 18630 24840
rect 18550 24660 18570 24820
rect 18610 24660 18630 24820
rect 18550 24640 18630 24660
rect 18660 24820 18740 24840
rect 18660 24660 18680 24820
rect 18720 24660 18740 24820
rect 18660 24640 18740 24660
rect 18770 24820 18850 24840
rect 18770 24660 18790 24820
rect 18830 24660 18850 24820
rect 18770 24640 18850 24660
rect 18880 24820 18960 24840
rect 18880 24660 18900 24820
rect 18940 24660 18960 24820
rect 18880 24640 18960 24660
rect 18990 24820 19070 24840
rect 18990 24660 19010 24820
rect 19050 24660 19070 24820
rect 18990 24640 19070 24660
rect 19100 24820 19180 24840
rect 19100 24660 19120 24820
rect 19160 24660 19180 24820
rect 19100 24640 19180 24660
rect 19210 24820 19290 24840
rect 19210 24660 19230 24820
rect 19270 24660 19290 24820
rect 19210 24640 19290 24660
rect 19320 24820 19400 24840
rect 19320 24660 19340 24820
rect 19380 24660 19400 24820
rect 19320 24640 19400 24660
rect 19430 24820 19510 24840
rect 19430 24660 19450 24820
rect 19490 24660 19510 24820
rect 19430 24640 19510 24660
rect 19540 24820 19620 24840
rect 19540 24660 19560 24820
rect 19600 24660 19620 24820
rect 19540 24640 19620 24660
rect 19650 24820 19730 24840
rect 19650 24660 19670 24820
rect 19710 24660 19730 24820
rect 19650 24640 19730 24660
rect 19760 24820 19840 24840
rect 19760 24660 19780 24820
rect 19820 24660 19840 24820
rect 19760 24640 19840 24660
rect 19870 24820 19950 24840
rect 19870 24660 19890 24820
rect 19930 24660 19950 24820
rect 19870 24640 19950 24660
rect 19980 24820 20060 24840
rect 19980 24660 20000 24820
rect 20040 24660 20060 24820
rect 19980 24640 20060 24660
rect 20090 24820 20170 24840
rect 20090 24660 20110 24820
rect 20150 24660 20170 24820
rect 20090 24640 20170 24660
rect 20200 24820 20280 24840
rect 20200 24660 20220 24820
rect 20260 24660 20280 24820
rect 20200 24640 20280 24660
rect 20310 24820 20390 24840
rect 20310 24660 20330 24820
rect 20370 24660 20390 24820
rect 20310 24640 20390 24660
rect 20420 24820 20500 24840
rect 20420 24660 20440 24820
rect 20480 24660 20500 24820
rect 20420 24640 20500 24660
rect 20530 24820 20600 24840
rect 20530 24660 20550 24820
rect 20590 24660 20600 24820
rect 20530 24640 20600 24660
rect 12150 24540 12220 24560
rect 12150 24380 12160 24540
rect 12200 24380 12220 24540
rect 12150 24360 12220 24380
rect 12250 24540 12330 24560
rect 12250 24380 12270 24540
rect 12310 24380 12330 24540
rect 12250 24360 12330 24380
rect 12360 24540 12430 24560
rect 12360 24380 12380 24540
rect 12420 24380 12430 24540
rect 12360 24360 12430 24380
rect 12530 24540 12600 24560
rect 12530 24380 12540 24540
rect 12580 24380 12600 24540
rect 12530 24360 12600 24380
rect 12630 24540 12710 24560
rect 12630 24380 12650 24540
rect 12690 24380 12710 24540
rect 12630 24360 12710 24380
rect 12740 24540 12810 24560
rect 12740 24380 12760 24540
rect 12800 24380 12810 24540
rect 12740 24360 12810 24380
rect 7360 22810 7430 23210
rect 7460 23190 7540 23210
rect 7460 22830 7480 23190
rect 7520 22830 7540 23190
rect 7460 22810 7540 22830
rect 7570 22810 7690 23210
rect 7720 23190 7800 23210
rect 7720 22830 7740 23190
rect 7780 22830 7800 23190
rect 7720 22810 7800 22830
rect 7830 22810 7900 23210
rect 7960 23190 8030 23210
rect 7960 23030 7970 23190
rect 8010 23030 8030 23190
rect 7960 23010 8030 23030
rect 8060 23190 8140 23210
rect 8060 23030 8080 23190
rect 8120 23030 8140 23190
rect 8060 23010 8140 23030
rect 8170 23190 8240 23210
rect 8170 23030 8190 23190
rect 8230 23030 8240 23190
rect 8170 23010 8240 23030
rect 8480 23190 8550 23210
rect 8480 22830 8490 23190
rect 8530 22830 8550 23190
rect 8480 22810 8550 22830
rect 8580 23190 8700 23210
rect 8580 22830 8620 23190
rect 8660 22830 8700 23190
rect 8580 22810 8700 22830
rect 8730 23190 8800 23210
rect 8730 22830 8750 23190
rect 8790 22830 8800 23190
rect 9220 23190 9290 23210
rect 9220 23030 9230 23190
rect 9270 23030 9290 23190
rect 9220 23010 9290 23030
rect 9320 23190 9400 23210
rect 9320 23030 9340 23190
rect 9380 23030 9400 23190
rect 9320 23010 9400 23030
rect 9430 23190 9500 23210
rect 9430 23030 9450 23190
rect 9490 23030 9500 23190
rect 9430 23010 9500 23030
rect 8730 22810 8800 22830
rect 8860 22920 8930 22940
rect 8860 22760 8870 22920
rect 8910 22760 8930 22920
rect 8860 22740 8930 22760
rect 8960 22920 9030 22940
rect 8960 22760 8980 22920
rect 9020 22760 9030 22920
rect 8960 22740 9030 22760
rect 9560 22810 9630 23210
rect 9660 23190 9740 23210
rect 9660 22830 9680 23190
rect 9720 22830 9740 23190
rect 9660 22810 9740 22830
rect 9770 22810 9890 23210
rect 9920 23190 10000 23210
rect 9920 22830 9940 23190
rect 9980 22830 10000 23190
rect 9920 22810 10000 22830
rect 10030 22810 10100 23210
rect 10160 23190 10230 23210
rect 10160 23030 10170 23190
rect 10210 23030 10230 23190
rect 10160 23010 10230 23030
rect 10260 23190 10340 23210
rect 10260 23030 10280 23190
rect 10320 23030 10340 23190
rect 10260 23010 10340 23030
rect 10370 23190 10440 23210
rect 10370 23030 10390 23190
rect 10430 23030 10440 23190
rect 10370 23010 10440 23030
rect 10550 22810 10620 23210
rect 10650 23190 10730 23210
rect 10650 22830 10670 23190
rect 10710 22830 10730 23190
rect 10650 22810 10730 22830
rect 10760 22810 10880 23210
rect 10910 23190 10990 23210
rect 10910 22830 10930 23190
rect 10970 22830 10990 23190
rect 10910 22810 10990 22830
rect 11020 22810 11090 23210
rect 11150 23190 11220 23210
rect 11150 23030 11160 23190
rect 11200 23030 11220 23190
rect 11150 23010 11220 23030
rect 11250 23190 11330 23210
rect 11250 23030 11270 23190
rect 11310 23030 11330 23190
rect 11250 23010 11330 23030
rect 11360 23190 11430 23210
rect 11360 23030 11380 23190
rect 11420 23030 11430 23190
rect 11360 23010 11430 23030
rect 11550 22810 11620 23210
rect 11650 23190 11730 23210
rect 11650 22830 11670 23190
rect 11710 22830 11730 23190
rect 11650 22810 11730 22830
rect 11760 22810 11880 23210
rect 11910 23190 11990 23210
rect 11910 22830 11930 23190
rect 11970 22830 11990 23190
rect 11910 22810 11990 22830
rect 12020 22810 12090 23210
rect 12150 23190 12220 23210
rect 12150 23030 12160 23190
rect 12200 23030 12220 23190
rect 12150 23010 12220 23030
rect 12250 23190 12330 23210
rect 12250 23030 12270 23190
rect 12310 23030 12330 23190
rect 12250 23010 12330 23030
rect 12360 23190 12430 23210
rect 12360 23030 12380 23190
rect 12420 23030 12430 23190
rect 12360 23010 12430 23030
rect 12530 23190 12600 23210
rect 12530 23030 12540 23190
rect 12580 23030 12600 23190
rect 12530 23010 12600 23030
rect 12630 23190 12710 23210
rect 12630 23030 12650 23190
rect 12690 23030 12710 23190
rect 12630 23010 12710 23030
rect 12740 23190 12810 23210
rect 12740 23030 12760 23190
rect 12800 23030 12810 23190
rect 12740 23010 12810 23030
rect 12880 22910 12950 22930
rect 12880 22750 12890 22910
rect 12930 22750 12950 22910
rect 12880 22730 12950 22750
rect 12980 22910 13050 22930
rect 12980 22750 13000 22910
rect 13040 22750 13050 22910
rect 12980 22730 13050 22750
rect 13110 22910 13180 22930
rect 13110 22750 13120 22910
rect 13160 22750 13180 22910
rect 13110 22730 13180 22750
rect 13210 22910 13290 22930
rect 13210 22750 13230 22910
rect 13270 22750 13290 22910
rect 13210 22730 13290 22750
rect 13320 22910 13390 22930
rect 13320 22750 13340 22910
rect 13380 22750 13390 22910
rect 13320 22730 13390 22750
rect 13450 22910 13520 22930
rect 13450 22750 13460 22910
rect 13500 22750 13520 22910
rect 13450 22730 13520 22750
rect 13550 22910 13630 22930
rect 13550 22750 13570 22910
rect 13610 22750 13630 22910
rect 13550 22730 13630 22750
rect 13660 22910 13740 22930
rect 13660 22750 13680 22910
rect 13720 22750 13740 22910
rect 13660 22730 13740 22750
rect 13770 22910 13850 22930
rect 13770 22750 13790 22910
rect 13830 22750 13850 22910
rect 13770 22730 13850 22750
rect 13880 22910 13950 22930
rect 13880 22750 13900 22910
rect 13940 22750 13950 22910
rect 13880 22730 13950 22750
rect 14010 22910 14080 22930
rect 14010 22750 14020 22910
rect 14060 22750 14080 22910
rect 14010 22730 14080 22750
rect 14110 22910 14190 22930
rect 14110 22750 14130 22910
rect 14170 22750 14190 22910
rect 14110 22730 14190 22750
rect 14220 22910 14300 22930
rect 14220 22750 14240 22910
rect 14280 22750 14300 22910
rect 14220 22730 14300 22750
rect 14330 22910 14410 22930
rect 14330 22750 14350 22910
rect 14390 22750 14410 22910
rect 14330 22730 14410 22750
rect 14440 22910 14520 22930
rect 14440 22750 14460 22910
rect 14500 22750 14520 22910
rect 14440 22730 14520 22750
rect 14550 22910 14630 22930
rect 14550 22750 14570 22910
rect 14610 22750 14630 22910
rect 14550 22730 14630 22750
rect 14660 22910 14740 22930
rect 14660 22750 14680 22910
rect 14720 22750 14740 22910
rect 14660 22730 14740 22750
rect 14770 22910 14850 22930
rect 14770 22750 14790 22910
rect 14830 22750 14850 22910
rect 14770 22730 14850 22750
rect 14880 22910 14950 22930
rect 14880 22750 14900 22910
rect 14940 22750 14950 22910
rect 14880 22730 14950 22750
rect 15070 22910 15140 22930
rect 15070 22750 15080 22910
rect 15120 22750 15140 22910
rect 15070 22730 15140 22750
rect 15170 22910 15250 22930
rect 15170 22750 15190 22910
rect 15230 22750 15250 22910
rect 15170 22730 15250 22750
rect 15280 22910 15360 22930
rect 15280 22750 15300 22910
rect 15340 22750 15360 22910
rect 15280 22730 15360 22750
rect 15390 22910 15470 22930
rect 15390 22750 15410 22910
rect 15450 22750 15470 22910
rect 15390 22730 15470 22750
rect 15500 22910 15580 22930
rect 15500 22750 15520 22910
rect 15560 22750 15580 22910
rect 15500 22730 15580 22750
rect 15610 22910 15690 22930
rect 15610 22750 15630 22910
rect 15670 22750 15690 22910
rect 15610 22730 15690 22750
rect 15720 22910 15800 22930
rect 15720 22750 15740 22910
rect 15780 22750 15800 22910
rect 15720 22730 15800 22750
rect 15830 22910 15910 22930
rect 15830 22750 15850 22910
rect 15890 22750 15910 22910
rect 15830 22730 15910 22750
rect 15940 22910 16020 22930
rect 15940 22750 15960 22910
rect 16000 22750 16020 22910
rect 15940 22730 16020 22750
rect 16050 22910 16130 22930
rect 16050 22750 16070 22910
rect 16110 22750 16130 22910
rect 16050 22730 16130 22750
rect 16160 22910 16240 22930
rect 16160 22750 16180 22910
rect 16220 22750 16240 22910
rect 16160 22730 16240 22750
rect 16270 22910 16350 22930
rect 16270 22750 16290 22910
rect 16330 22750 16350 22910
rect 16270 22730 16350 22750
rect 16380 22910 16460 22930
rect 16380 22750 16400 22910
rect 16440 22750 16460 22910
rect 16380 22730 16460 22750
rect 16490 22910 16570 22930
rect 16490 22750 16510 22910
rect 16550 22750 16570 22910
rect 16490 22730 16570 22750
rect 16600 22910 16680 22930
rect 16600 22750 16620 22910
rect 16660 22750 16680 22910
rect 16600 22730 16680 22750
rect 16710 22910 16790 22930
rect 16710 22750 16730 22910
rect 16770 22750 16790 22910
rect 16710 22730 16790 22750
rect 16820 22910 16890 22930
rect 16820 22750 16840 22910
rect 16880 22750 16890 22910
rect 16820 22730 16890 22750
rect 17020 22910 17090 22930
rect 17020 22750 17030 22910
rect 17070 22750 17090 22910
rect 17020 22730 17090 22750
rect 17120 22910 17200 22930
rect 17120 22750 17140 22910
rect 17180 22750 17200 22910
rect 17120 22730 17200 22750
rect 17230 22910 17310 22930
rect 17230 22750 17250 22910
rect 17290 22750 17310 22910
rect 17230 22730 17310 22750
rect 17340 22910 17420 22930
rect 17340 22750 17360 22910
rect 17400 22750 17420 22910
rect 17340 22730 17420 22750
rect 17450 22910 17530 22930
rect 17450 22750 17470 22910
rect 17510 22750 17530 22910
rect 17450 22730 17530 22750
rect 17560 22910 17640 22930
rect 17560 22750 17580 22910
rect 17620 22750 17640 22910
rect 17560 22730 17640 22750
rect 17670 22910 17750 22930
rect 17670 22750 17690 22910
rect 17730 22750 17750 22910
rect 17670 22730 17750 22750
rect 17780 22910 17860 22930
rect 17780 22750 17800 22910
rect 17840 22750 17860 22910
rect 17780 22730 17860 22750
rect 17890 22910 17970 22930
rect 17890 22750 17910 22910
rect 17950 22750 17970 22910
rect 17890 22730 17970 22750
rect 18000 22910 18080 22930
rect 18000 22750 18020 22910
rect 18060 22750 18080 22910
rect 18000 22730 18080 22750
rect 18110 22910 18190 22930
rect 18110 22750 18130 22910
rect 18170 22750 18190 22910
rect 18110 22730 18190 22750
rect 18220 22910 18300 22930
rect 18220 22750 18240 22910
rect 18280 22750 18300 22910
rect 18220 22730 18300 22750
rect 18330 22910 18410 22930
rect 18330 22750 18350 22910
rect 18390 22750 18410 22910
rect 18330 22730 18410 22750
rect 18440 22910 18520 22930
rect 18440 22750 18460 22910
rect 18500 22750 18520 22910
rect 18440 22730 18520 22750
rect 18550 22910 18630 22930
rect 18550 22750 18570 22910
rect 18610 22750 18630 22910
rect 18550 22730 18630 22750
rect 18660 22910 18740 22930
rect 18660 22750 18680 22910
rect 18720 22750 18740 22910
rect 18660 22730 18740 22750
rect 18770 22910 18850 22930
rect 18770 22750 18790 22910
rect 18830 22750 18850 22910
rect 18770 22730 18850 22750
rect 18880 22910 18960 22930
rect 18880 22750 18900 22910
rect 18940 22750 18960 22910
rect 18880 22730 18960 22750
rect 18990 22910 19070 22930
rect 18990 22750 19010 22910
rect 19050 22750 19070 22910
rect 18990 22730 19070 22750
rect 19100 22910 19180 22930
rect 19100 22750 19120 22910
rect 19160 22750 19180 22910
rect 19100 22730 19180 22750
rect 19210 22910 19290 22930
rect 19210 22750 19230 22910
rect 19270 22750 19290 22910
rect 19210 22730 19290 22750
rect 19320 22910 19400 22930
rect 19320 22750 19340 22910
rect 19380 22750 19400 22910
rect 19320 22730 19400 22750
rect 19430 22910 19510 22930
rect 19430 22750 19450 22910
rect 19490 22750 19510 22910
rect 19430 22730 19510 22750
rect 19540 22910 19620 22930
rect 19540 22750 19560 22910
rect 19600 22750 19620 22910
rect 19540 22730 19620 22750
rect 19650 22910 19730 22930
rect 19650 22750 19670 22910
rect 19710 22750 19730 22910
rect 19650 22730 19730 22750
rect 19760 22910 19840 22930
rect 19760 22750 19780 22910
rect 19820 22750 19840 22910
rect 19760 22730 19840 22750
rect 19870 22910 19950 22930
rect 19870 22750 19890 22910
rect 19930 22750 19950 22910
rect 19870 22730 19950 22750
rect 19980 22910 20060 22930
rect 19980 22750 20000 22910
rect 20040 22750 20060 22910
rect 19980 22730 20060 22750
rect 20090 22910 20170 22930
rect 20090 22750 20110 22910
rect 20150 22750 20170 22910
rect 20090 22730 20170 22750
rect 20200 22910 20280 22930
rect 20200 22750 20220 22910
rect 20260 22750 20280 22910
rect 20200 22730 20280 22750
rect 20310 22910 20390 22930
rect 20310 22750 20330 22910
rect 20370 22750 20390 22910
rect 20310 22730 20390 22750
rect 20420 22910 20500 22930
rect 20420 22750 20440 22910
rect 20480 22750 20500 22910
rect 20420 22730 20500 22750
rect 20530 22910 20600 22930
rect 20530 22750 20550 22910
rect 20590 22750 20600 22910
rect 20530 22730 20600 22750
rect 8860 18220 8930 18240
rect 8480 18150 8550 18170
rect 7280 17960 7350 17980
rect 7280 17800 7290 17960
rect 7330 17800 7350 17960
rect 7280 17780 7350 17800
rect 7380 17960 7460 17980
rect 7380 17800 7400 17960
rect 7440 17800 7460 17960
rect 7380 17780 7460 17800
rect 7490 17960 7610 17980
rect 7490 17800 7530 17960
rect 7570 17800 7610 17960
rect 7490 17780 7610 17800
rect 7640 17960 7720 17980
rect 7640 17800 7660 17960
rect 7700 17800 7720 17960
rect 7640 17780 7720 17800
rect 7750 17960 7820 17980
rect 7750 17800 7770 17960
rect 7810 17800 7820 17960
rect 7750 17780 7820 17800
rect 7950 17960 8020 17980
rect 7950 17800 7960 17960
rect 8000 17800 8020 17960
rect 7950 17780 8020 17800
rect 8050 17960 8130 17980
rect 8050 17800 8070 17960
rect 8110 17800 8130 17960
rect 8050 17780 8130 17800
rect 8160 17960 8230 17980
rect 8160 17800 8180 17960
rect 8220 17800 8230 17960
rect 8160 17780 8230 17800
rect 8480 17790 8490 18150
rect 8530 17790 8550 18150
rect 8480 17770 8550 17790
rect 8580 18150 8700 18170
rect 8580 17790 8620 18150
rect 8660 17790 8700 18150
rect 8580 17770 8700 17790
rect 8730 18150 8800 18170
rect 8730 17790 8750 18150
rect 8790 17790 8800 18150
rect 8860 18060 8870 18220
rect 8910 18060 8930 18220
rect 8860 18040 8930 18060
rect 8960 18220 9030 18240
rect 8960 18060 8980 18220
rect 9020 18060 9030 18220
rect 8960 18040 9030 18060
rect 8730 17770 8800 17790
rect 9220 17950 9290 17970
rect 9220 17790 9230 17950
rect 9270 17790 9290 17950
rect 9220 17770 9290 17790
rect 9320 17950 9400 17970
rect 9320 17790 9340 17950
rect 9380 17790 9400 17950
rect 9320 17770 9400 17790
rect 9430 17950 9500 17970
rect 9430 17790 9450 17950
rect 9490 17790 9500 17950
rect 9430 17770 9500 17790
rect 9560 17770 9630 18170
rect 9660 18150 9740 18170
rect 9660 17790 9680 18150
rect 9720 17790 9740 18150
rect 9660 17770 9740 17790
rect 9770 17770 9890 18170
rect 9920 18150 10000 18170
rect 9920 17790 9940 18150
rect 9980 17790 10000 18150
rect 9920 17770 10000 17790
rect 10030 17770 10100 18170
rect 10160 17950 10230 17970
rect 10160 17790 10170 17950
rect 10210 17790 10230 17950
rect 10160 17770 10230 17790
rect 10260 17950 10340 17970
rect 10260 17790 10280 17950
rect 10320 17790 10340 17950
rect 10260 17770 10340 17790
rect 10370 17950 10440 17970
rect 10370 17790 10390 17950
rect 10430 17790 10440 17950
rect 10370 17770 10440 17790
rect 10550 17770 10620 18170
rect 10650 18150 10730 18170
rect 10650 17790 10670 18150
rect 10710 17790 10730 18150
rect 10650 17770 10730 17790
rect 10760 17770 10880 18170
rect 10910 18150 10990 18170
rect 10910 17790 10930 18150
rect 10970 17790 10990 18150
rect 10910 17770 10990 17790
rect 11020 17770 11090 18170
rect 11150 17950 11220 17970
rect 11150 17790 11160 17950
rect 11200 17790 11220 17950
rect 11150 17770 11220 17790
rect 11250 17950 11330 17970
rect 11250 17790 11270 17950
rect 11310 17790 11330 17950
rect 11250 17770 11330 17790
rect 11360 17950 11430 17970
rect 11360 17790 11380 17950
rect 11420 17790 11430 17950
rect 11360 17770 11430 17790
rect 11550 17770 11620 18170
rect 11650 18150 11730 18170
rect 11650 17790 11670 18150
rect 11710 17790 11730 18150
rect 11650 17770 11730 17790
rect 11760 17770 11880 18170
rect 11910 18150 11990 18170
rect 11910 17790 11930 18150
rect 11970 17790 11990 18150
rect 11910 17770 11990 17790
rect 12020 17770 12090 18170
rect 12880 18230 12950 18250
rect 12880 18070 12890 18230
rect 12930 18070 12950 18230
rect 12880 18050 12950 18070
rect 12980 18230 13050 18250
rect 12980 18070 13000 18230
rect 13040 18070 13050 18230
rect 12980 18050 13050 18070
rect 13110 18230 13180 18250
rect 13110 18070 13120 18230
rect 13160 18070 13180 18230
rect 13110 18050 13180 18070
rect 13210 18230 13290 18250
rect 13210 18070 13230 18230
rect 13270 18070 13290 18230
rect 13210 18050 13290 18070
rect 13320 18230 13390 18250
rect 13320 18070 13340 18230
rect 13380 18070 13390 18230
rect 13320 18050 13390 18070
rect 13450 18230 13520 18250
rect 13450 18070 13460 18230
rect 13500 18070 13520 18230
rect 13450 18050 13520 18070
rect 13550 18230 13630 18250
rect 13550 18070 13570 18230
rect 13610 18070 13630 18230
rect 13550 18050 13630 18070
rect 13660 18230 13740 18250
rect 13660 18070 13680 18230
rect 13720 18070 13740 18230
rect 13660 18050 13740 18070
rect 13770 18230 13850 18250
rect 13770 18070 13790 18230
rect 13830 18070 13850 18230
rect 13770 18050 13850 18070
rect 13880 18230 13950 18250
rect 13880 18070 13900 18230
rect 13940 18070 13950 18230
rect 13880 18050 13950 18070
rect 14010 18230 14080 18250
rect 14010 18070 14020 18230
rect 14060 18070 14080 18230
rect 14010 18050 14080 18070
rect 14110 18230 14190 18250
rect 14110 18070 14130 18230
rect 14170 18070 14190 18230
rect 14110 18050 14190 18070
rect 14220 18230 14300 18250
rect 14220 18070 14240 18230
rect 14280 18070 14300 18230
rect 14220 18050 14300 18070
rect 14330 18230 14410 18250
rect 14330 18070 14350 18230
rect 14390 18070 14410 18230
rect 14330 18050 14410 18070
rect 14440 18230 14520 18250
rect 14440 18070 14460 18230
rect 14500 18070 14520 18230
rect 14440 18050 14520 18070
rect 14550 18230 14630 18250
rect 14550 18070 14570 18230
rect 14610 18070 14630 18230
rect 14550 18050 14630 18070
rect 14660 18230 14740 18250
rect 14660 18070 14680 18230
rect 14720 18070 14740 18230
rect 14660 18050 14740 18070
rect 14770 18230 14850 18250
rect 14770 18070 14790 18230
rect 14830 18070 14850 18230
rect 14770 18050 14850 18070
rect 14880 18230 14950 18250
rect 14880 18070 14900 18230
rect 14940 18070 14950 18230
rect 14880 18050 14950 18070
rect 15070 18230 15140 18250
rect 15070 18070 15080 18230
rect 15120 18070 15140 18230
rect 15070 18050 15140 18070
rect 15170 18230 15250 18250
rect 15170 18070 15190 18230
rect 15230 18070 15250 18230
rect 15170 18050 15250 18070
rect 15280 18230 15360 18250
rect 15280 18070 15300 18230
rect 15340 18070 15360 18230
rect 15280 18050 15360 18070
rect 15390 18230 15470 18250
rect 15390 18070 15410 18230
rect 15450 18070 15470 18230
rect 15390 18050 15470 18070
rect 15500 18230 15580 18250
rect 15500 18070 15520 18230
rect 15560 18070 15580 18230
rect 15500 18050 15580 18070
rect 15610 18230 15690 18250
rect 15610 18070 15630 18230
rect 15670 18070 15690 18230
rect 15610 18050 15690 18070
rect 15720 18230 15800 18250
rect 15720 18070 15740 18230
rect 15780 18070 15800 18230
rect 15720 18050 15800 18070
rect 15830 18230 15910 18250
rect 15830 18070 15850 18230
rect 15890 18070 15910 18230
rect 15830 18050 15910 18070
rect 15940 18230 16020 18250
rect 15940 18070 15960 18230
rect 16000 18070 16020 18230
rect 15940 18050 16020 18070
rect 16050 18230 16130 18250
rect 16050 18070 16070 18230
rect 16110 18070 16130 18230
rect 16050 18050 16130 18070
rect 16160 18230 16240 18250
rect 16160 18070 16180 18230
rect 16220 18070 16240 18230
rect 16160 18050 16240 18070
rect 16270 18230 16350 18250
rect 16270 18070 16290 18230
rect 16330 18070 16350 18230
rect 16270 18050 16350 18070
rect 16380 18230 16460 18250
rect 16380 18070 16400 18230
rect 16440 18070 16460 18230
rect 16380 18050 16460 18070
rect 16490 18230 16570 18250
rect 16490 18070 16510 18230
rect 16550 18070 16570 18230
rect 16490 18050 16570 18070
rect 16600 18230 16680 18250
rect 16600 18070 16620 18230
rect 16660 18070 16680 18230
rect 16600 18050 16680 18070
rect 16710 18230 16790 18250
rect 16710 18070 16730 18230
rect 16770 18070 16790 18230
rect 16710 18050 16790 18070
rect 16820 18230 16890 18250
rect 16820 18070 16840 18230
rect 16880 18070 16890 18230
rect 16820 18050 16890 18070
rect 17020 18230 17090 18250
rect 17020 18070 17030 18230
rect 17070 18070 17090 18230
rect 17020 18050 17090 18070
rect 17120 18230 17200 18250
rect 17120 18070 17140 18230
rect 17180 18070 17200 18230
rect 17120 18050 17200 18070
rect 17230 18230 17310 18250
rect 17230 18070 17250 18230
rect 17290 18070 17310 18230
rect 17230 18050 17310 18070
rect 17340 18230 17420 18250
rect 17340 18070 17360 18230
rect 17400 18070 17420 18230
rect 17340 18050 17420 18070
rect 17450 18230 17530 18250
rect 17450 18070 17470 18230
rect 17510 18070 17530 18230
rect 17450 18050 17530 18070
rect 17560 18230 17640 18250
rect 17560 18070 17580 18230
rect 17620 18070 17640 18230
rect 17560 18050 17640 18070
rect 17670 18230 17750 18250
rect 17670 18070 17690 18230
rect 17730 18070 17750 18230
rect 17670 18050 17750 18070
rect 17780 18230 17860 18250
rect 17780 18070 17800 18230
rect 17840 18070 17860 18230
rect 17780 18050 17860 18070
rect 17890 18230 17970 18250
rect 17890 18070 17910 18230
rect 17950 18070 17970 18230
rect 17890 18050 17970 18070
rect 18000 18230 18080 18250
rect 18000 18070 18020 18230
rect 18060 18070 18080 18230
rect 18000 18050 18080 18070
rect 18110 18230 18190 18250
rect 18110 18070 18130 18230
rect 18170 18070 18190 18230
rect 18110 18050 18190 18070
rect 18220 18230 18300 18250
rect 18220 18070 18240 18230
rect 18280 18070 18300 18230
rect 18220 18050 18300 18070
rect 18330 18230 18410 18250
rect 18330 18070 18350 18230
rect 18390 18070 18410 18230
rect 18330 18050 18410 18070
rect 18440 18230 18520 18250
rect 18440 18070 18460 18230
rect 18500 18070 18520 18230
rect 18440 18050 18520 18070
rect 18550 18230 18630 18250
rect 18550 18070 18570 18230
rect 18610 18070 18630 18230
rect 18550 18050 18630 18070
rect 18660 18230 18740 18250
rect 18660 18070 18680 18230
rect 18720 18070 18740 18230
rect 18660 18050 18740 18070
rect 18770 18230 18850 18250
rect 18770 18070 18790 18230
rect 18830 18070 18850 18230
rect 18770 18050 18850 18070
rect 18880 18230 18960 18250
rect 18880 18070 18900 18230
rect 18940 18070 18960 18230
rect 18880 18050 18960 18070
rect 18990 18230 19070 18250
rect 18990 18070 19010 18230
rect 19050 18070 19070 18230
rect 18990 18050 19070 18070
rect 19100 18230 19180 18250
rect 19100 18070 19120 18230
rect 19160 18070 19180 18230
rect 19100 18050 19180 18070
rect 19210 18230 19290 18250
rect 19210 18070 19230 18230
rect 19270 18070 19290 18230
rect 19210 18050 19290 18070
rect 19320 18230 19400 18250
rect 19320 18070 19340 18230
rect 19380 18070 19400 18230
rect 19320 18050 19400 18070
rect 19430 18230 19510 18250
rect 19430 18070 19450 18230
rect 19490 18070 19510 18230
rect 19430 18050 19510 18070
rect 19540 18230 19620 18250
rect 19540 18070 19560 18230
rect 19600 18070 19620 18230
rect 19540 18050 19620 18070
rect 19650 18230 19730 18250
rect 19650 18070 19670 18230
rect 19710 18070 19730 18230
rect 19650 18050 19730 18070
rect 19760 18230 19840 18250
rect 19760 18070 19780 18230
rect 19820 18070 19840 18230
rect 19760 18050 19840 18070
rect 19870 18230 19950 18250
rect 19870 18070 19890 18230
rect 19930 18070 19950 18230
rect 19870 18050 19950 18070
rect 19980 18230 20060 18250
rect 19980 18070 20000 18230
rect 20040 18070 20060 18230
rect 19980 18050 20060 18070
rect 20090 18230 20170 18250
rect 20090 18070 20110 18230
rect 20150 18070 20170 18230
rect 20090 18050 20170 18070
rect 20200 18230 20280 18250
rect 20200 18070 20220 18230
rect 20260 18070 20280 18230
rect 20200 18050 20280 18070
rect 20310 18230 20390 18250
rect 20310 18070 20330 18230
rect 20370 18070 20390 18230
rect 20310 18050 20390 18070
rect 20420 18230 20500 18250
rect 20420 18070 20440 18230
rect 20480 18070 20500 18230
rect 20420 18050 20500 18070
rect 20530 18230 20600 18250
rect 20530 18070 20550 18230
rect 20590 18070 20600 18230
rect 20530 18050 20600 18070
rect 12150 17950 12220 17970
rect 12150 17790 12160 17950
rect 12200 17790 12220 17950
rect 12150 17770 12220 17790
rect 12250 17950 12330 17970
rect 12250 17790 12270 17950
rect 12310 17790 12330 17950
rect 12250 17770 12330 17790
rect 12360 17950 12430 17970
rect 12360 17790 12380 17950
rect 12420 17790 12430 17950
rect 12360 17770 12430 17790
rect 12530 17950 12600 17970
rect 12530 17790 12540 17950
rect 12580 17790 12600 17950
rect 12530 17770 12600 17790
rect 12630 17950 12710 17970
rect 12630 17790 12650 17950
rect 12690 17790 12710 17950
rect 12630 17770 12710 17790
rect 12740 17950 12810 17970
rect 12740 17790 12760 17950
rect 12800 17790 12810 17950
rect 12740 17770 12810 17790
rect 9760 15530 9830 15550
rect 9760 15370 9770 15530
rect 9810 15370 9830 15530
rect 9760 15350 9830 15370
rect 9860 15530 9940 15550
rect 9860 15370 9880 15530
rect 9920 15370 9940 15530
rect 9860 15350 9940 15370
rect 9970 15530 10040 15550
rect 9970 15370 9990 15530
rect 10030 15370 10040 15530
rect 9970 15350 10040 15370
rect 10300 15150 10370 15550
rect 10400 15530 10480 15550
rect 10400 15170 10420 15530
rect 10460 15170 10480 15530
rect 10400 15150 10480 15170
rect 10510 15150 10630 15550
rect 10660 15530 10740 15550
rect 10660 15170 10680 15530
rect 10720 15170 10740 15530
rect 10660 15150 10740 15170
rect 10770 15150 10840 15550
rect 10900 15530 10970 15550
rect 10900 15370 10910 15530
rect 10950 15370 10970 15530
rect 10900 15350 10970 15370
rect 11000 15530 11080 15550
rect 11000 15370 11020 15530
rect 11060 15370 11080 15530
rect 11000 15350 11080 15370
rect 11110 15530 11180 15550
rect 11110 15370 11130 15530
rect 11170 15370 11180 15530
rect 11110 15350 11180 15370
rect 11290 15150 11360 15550
rect 11390 15530 11470 15550
rect 11390 15170 11410 15530
rect 11450 15170 11470 15530
rect 11390 15150 11470 15170
rect 11500 15150 11620 15550
rect 11650 15530 11730 15550
rect 11650 15170 11670 15530
rect 11710 15170 11730 15530
rect 11650 15150 11730 15170
rect 11760 15150 11830 15550
rect 11890 15530 11960 15550
rect 11890 15370 11900 15530
rect 11940 15370 11960 15530
rect 11890 15350 11960 15370
rect 11990 15530 12070 15550
rect 11990 15370 12010 15530
rect 12050 15370 12070 15530
rect 11990 15350 12070 15370
rect 12100 15530 12170 15550
rect 12100 15370 12120 15530
rect 12160 15370 12170 15530
rect 12100 15350 12170 15370
rect 12290 15150 12360 15550
rect 12390 15530 12470 15550
rect 12390 15170 12410 15530
rect 12450 15170 12470 15530
rect 12390 15150 12470 15170
rect 12500 15150 12620 15550
rect 12650 15530 12730 15550
rect 12650 15170 12670 15530
rect 12710 15170 12730 15530
rect 12650 15150 12730 15170
rect 12760 15150 12830 15550
rect 12890 15530 12960 15550
rect 12890 15370 12900 15530
rect 12940 15370 12960 15530
rect 12890 15350 12960 15370
rect 12990 15530 13070 15550
rect 12990 15370 13010 15530
rect 13050 15370 13070 15530
rect 12990 15350 13070 15370
rect 13100 15530 13170 15550
rect 13100 15370 13120 15530
rect 13160 15370 13170 15530
rect 13100 15350 13170 15370
rect 13240 15250 13310 15270
rect 13240 15090 13250 15250
rect 13290 15090 13310 15250
rect 13240 15070 13310 15090
rect 13340 15250 13410 15270
rect 13340 15090 13360 15250
rect 13400 15090 13410 15250
rect 13340 15070 13410 15090
rect 13470 15250 13540 15270
rect 13470 15090 13480 15250
rect 13520 15090 13540 15250
rect 13470 15070 13540 15090
rect 13570 15250 13650 15270
rect 13570 15090 13590 15250
rect 13630 15090 13650 15250
rect 13570 15070 13650 15090
rect 13680 15250 13750 15270
rect 13680 15090 13700 15250
rect 13740 15090 13750 15250
rect 13680 15070 13750 15090
rect 13810 15250 13880 15270
rect 13810 15090 13820 15250
rect 13860 15090 13880 15250
rect 13810 15070 13880 15090
rect 13910 15250 13990 15270
rect 13910 15090 13930 15250
rect 13970 15090 13990 15250
rect 13910 15070 13990 15090
rect 14020 15250 14100 15270
rect 14020 15090 14040 15250
rect 14080 15090 14100 15250
rect 14020 15070 14100 15090
rect 14130 15250 14210 15270
rect 14130 15090 14150 15250
rect 14190 15090 14210 15250
rect 14130 15070 14210 15090
rect 14240 15250 14310 15270
rect 14240 15090 14260 15250
rect 14300 15090 14310 15250
rect 14240 15070 14310 15090
rect 14370 15250 14440 15270
rect 14370 15090 14380 15250
rect 14420 15090 14440 15250
rect 14370 15070 14440 15090
rect 14470 15250 14550 15270
rect 14470 15090 14490 15250
rect 14530 15090 14550 15250
rect 14470 15070 14550 15090
rect 14580 15250 14660 15270
rect 14580 15090 14600 15250
rect 14640 15090 14660 15250
rect 14580 15070 14660 15090
rect 14690 15250 14770 15270
rect 14690 15090 14710 15250
rect 14750 15090 14770 15250
rect 14690 15070 14770 15090
rect 14800 15250 14880 15270
rect 14800 15090 14820 15250
rect 14860 15090 14880 15250
rect 14800 15070 14880 15090
rect 14910 15250 14990 15270
rect 14910 15090 14930 15250
rect 14970 15090 14990 15250
rect 14910 15070 14990 15090
rect 15020 15250 15100 15270
rect 15020 15090 15040 15250
rect 15080 15090 15100 15250
rect 15020 15070 15100 15090
rect 15130 15250 15210 15270
rect 15130 15090 15150 15250
rect 15190 15090 15210 15250
rect 15130 15070 15210 15090
rect 15240 15250 15310 15270
rect 15240 15090 15260 15250
rect 15300 15090 15310 15250
rect 15240 15070 15310 15090
rect 15430 15250 15500 15270
rect 15430 15090 15440 15250
rect 15480 15090 15500 15250
rect 15430 15070 15500 15090
rect 15530 15250 15610 15270
rect 15530 15090 15550 15250
rect 15590 15090 15610 15250
rect 15530 15070 15610 15090
rect 15640 15250 15720 15270
rect 15640 15090 15660 15250
rect 15700 15090 15720 15250
rect 15640 15070 15720 15090
rect 15750 15250 15830 15270
rect 15750 15090 15770 15250
rect 15810 15090 15830 15250
rect 15750 15070 15830 15090
rect 15860 15250 15940 15270
rect 15860 15090 15880 15250
rect 15920 15090 15940 15250
rect 15860 15070 15940 15090
rect 15970 15250 16050 15270
rect 15970 15090 15990 15250
rect 16030 15090 16050 15250
rect 15970 15070 16050 15090
rect 16080 15250 16160 15270
rect 16080 15090 16100 15250
rect 16140 15090 16160 15250
rect 16080 15070 16160 15090
rect 16190 15250 16270 15270
rect 16190 15090 16210 15250
rect 16250 15090 16270 15250
rect 16190 15070 16270 15090
rect 16300 15250 16380 15270
rect 16300 15090 16320 15250
rect 16360 15090 16380 15250
rect 16300 15070 16380 15090
rect 16410 15250 16490 15270
rect 16410 15090 16430 15250
rect 16470 15090 16490 15250
rect 16410 15070 16490 15090
rect 16520 15250 16600 15270
rect 16520 15090 16540 15250
rect 16580 15090 16600 15250
rect 16520 15070 16600 15090
rect 16630 15250 16710 15270
rect 16630 15090 16650 15250
rect 16690 15090 16710 15250
rect 16630 15070 16710 15090
rect 16740 15250 16820 15270
rect 16740 15090 16760 15250
rect 16800 15090 16820 15250
rect 16740 15070 16820 15090
rect 16850 15250 16930 15270
rect 16850 15090 16870 15250
rect 16910 15090 16930 15250
rect 16850 15070 16930 15090
rect 16960 15250 17040 15270
rect 16960 15090 16980 15250
rect 17020 15090 17040 15250
rect 16960 15070 17040 15090
rect 17070 15250 17150 15270
rect 17070 15090 17090 15250
rect 17130 15090 17150 15250
rect 17070 15070 17150 15090
rect 17180 15250 17250 15270
rect 17180 15090 17200 15250
rect 17240 15090 17250 15250
rect 17180 15070 17250 15090
rect 17380 15250 17450 15270
rect 17380 15090 17390 15250
rect 17430 15090 17450 15250
rect 17380 15070 17450 15090
rect 17480 15250 17560 15270
rect 17480 15090 17500 15250
rect 17540 15090 17560 15250
rect 17480 15070 17560 15090
rect 17590 15250 17670 15270
rect 17590 15090 17610 15250
rect 17650 15090 17670 15250
rect 17590 15070 17670 15090
rect 17700 15250 17780 15270
rect 17700 15090 17720 15250
rect 17760 15090 17780 15250
rect 17700 15070 17780 15090
rect 17810 15250 17890 15270
rect 17810 15090 17830 15250
rect 17870 15090 17890 15250
rect 17810 15070 17890 15090
rect 17920 15250 18000 15270
rect 17920 15090 17940 15250
rect 17980 15090 18000 15250
rect 17920 15070 18000 15090
rect 18030 15250 18110 15270
rect 18030 15090 18050 15250
rect 18090 15090 18110 15250
rect 18030 15070 18110 15090
rect 18140 15250 18220 15270
rect 18140 15090 18160 15250
rect 18200 15090 18220 15250
rect 18140 15070 18220 15090
rect 18250 15250 18330 15270
rect 18250 15090 18270 15250
rect 18310 15090 18330 15250
rect 18250 15070 18330 15090
rect 18360 15250 18440 15270
rect 18360 15090 18380 15250
rect 18420 15090 18440 15250
rect 18360 15070 18440 15090
rect 18470 15250 18550 15270
rect 18470 15090 18490 15250
rect 18530 15090 18550 15250
rect 18470 15070 18550 15090
rect 18580 15250 18660 15270
rect 18580 15090 18600 15250
rect 18640 15090 18660 15250
rect 18580 15070 18660 15090
rect 18690 15250 18770 15270
rect 18690 15090 18710 15250
rect 18750 15090 18770 15250
rect 18690 15070 18770 15090
rect 18800 15250 18880 15270
rect 18800 15090 18820 15250
rect 18860 15090 18880 15250
rect 18800 15070 18880 15090
rect 18910 15250 18990 15270
rect 18910 15090 18930 15250
rect 18970 15090 18990 15250
rect 18910 15070 18990 15090
rect 19020 15250 19100 15270
rect 19020 15090 19040 15250
rect 19080 15090 19100 15250
rect 19020 15070 19100 15090
rect 19130 15250 19210 15270
rect 19130 15090 19150 15250
rect 19190 15090 19210 15250
rect 19130 15070 19210 15090
rect 19240 15250 19320 15270
rect 19240 15090 19260 15250
rect 19300 15090 19320 15250
rect 19240 15070 19320 15090
rect 19350 15250 19430 15270
rect 19350 15090 19370 15250
rect 19410 15090 19430 15250
rect 19350 15070 19430 15090
rect 19460 15250 19540 15270
rect 19460 15090 19480 15250
rect 19520 15090 19540 15250
rect 19460 15070 19540 15090
rect 19570 15250 19650 15270
rect 19570 15090 19590 15250
rect 19630 15090 19650 15250
rect 19570 15070 19650 15090
rect 19680 15250 19760 15270
rect 19680 15090 19700 15250
rect 19740 15090 19760 15250
rect 19680 15070 19760 15090
rect 19790 15250 19870 15270
rect 19790 15090 19810 15250
rect 19850 15090 19870 15250
rect 19790 15070 19870 15090
rect 19900 15250 19980 15270
rect 19900 15090 19920 15250
rect 19960 15090 19980 15250
rect 19900 15070 19980 15090
rect 20010 15250 20090 15270
rect 20010 15090 20030 15250
rect 20070 15090 20090 15250
rect 20010 15070 20090 15090
rect 20120 15250 20200 15270
rect 20120 15090 20140 15250
rect 20180 15090 20200 15250
rect 20120 15070 20200 15090
rect 20230 15250 20310 15270
rect 20230 15090 20250 15250
rect 20290 15090 20310 15250
rect 20230 15070 20310 15090
rect 20340 15250 20420 15270
rect 20340 15090 20360 15250
rect 20400 15090 20420 15250
rect 20340 15070 20420 15090
rect 20450 15250 20530 15270
rect 20450 15090 20470 15250
rect 20510 15090 20530 15250
rect 20450 15070 20530 15090
rect 20560 15250 20640 15270
rect 20560 15090 20580 15250
rect 20620 15090 20640 15250
rect 20560 15070 20640 15090
rect 20670 15250 20750 15270
rect 20670 15090 20690 15250
rect 20730 15090 20750 15250
rect 20670 15070 20750 15090
rect 20780 15250 20860 15270
rect 20780 15090 20800 15250
rect 20840 15090 20860 15250
rect 20780 15070 20860 15090
rect 20890 15250 20960 15270
rect 20890 15090 20910 15250
rect 20950 15090 20960 15250
rect 20890 15070 20960 15090
rect 7280 12300 7350 12320
rect 7280 12140 7290 12300
rect 7330 12140 7350 12300
rect 7280 12120 7350 12140
rect 7380 12300 7460 12320
rect 7380 12140 7400 12300
rect 7440 12140 7460 12300
rect 7380 12120 7460 12140
rect 7490 12300 7560 12320
rect 7490 12140 7510 12300
rect 7550 12140 7560 12300
rect 7490 12120 7560 12140
rect 7800 12120 7870 12520
rect 7900 12500 7980 12520
rect 7900 12140 7920 12500
rect 7960 12140 7980 12500
rect 7900 12120 7980 12140
rect 8010 12120 8130 12520
rect 8160 12500 8240 12520
rect 8160 12140 8180 12500
rect 8220 12140 8240 12500
rect 8160 12120 8240 12140
rect 8270 12120 8340 12520
rect 8930 12570 9000 12590
rect 8550 12460 8620 12480
rect 8550 12100 8560 12460
rect 8600 12100 8620 12460
rect 8550 12080 8620 12100
rect 8650 12460 8770 12480
rect 8650 12100 8690 12460
rect 8730 12100 8770 12460
rect 8650 12080 8770 12100
rect 8800 12460 8870 12480
rect 8800 12100 8820 12460
rect 8860 12100 8870 12460
rect 8930 12410 8940 12570
rect 8980 12410 9000 12570
rect 8930 12390 9000 12410
rect 9030 12570 9100 12590
rect 9030 12410 9050 12570
rect 9090 12410 9100 12570
rect 9030 12390 9100 12410
rect 9190 12570 9260 12590
rect 9190 12410 9200 12570
rect 9240 12410 9260 12570
rect 9190 12390 9260 12410
rect 9290 12570 9360 12590
rect 9290 12410 9310 12570
rect 9350 12410 9360 12570
rect 9290 12390 9360 12410
rect 9440 12570 9510 12590
rect 9440 12410 9450 12570
rect 9490 12410 9510 12570
rect 9440 12390 9510 12410
rect 9540 12570 9610 12590
rect 9540 12410 9560 12570
rect 9600 12410 9610 12570
rect 9540 12390 9610 12410
rect 9860 12300 9930 12320
rect 9860 12140 9870 12300
rect 9910 12140 9930 12300
rect 9860 12120 9930 12140
rect 9960 12300 10040 12320
rect 9960 12140 9980 12300
rect 10020 12140 10040 12300
rect 9960 12120 10040 12140
rect 10070 12300 10140 12320
rect 10070 12140 10090 12300
rect 10130 12140 10140 12300
rect 10070 12120 10140 12140
rect 10400 12120 10470 12520
rect 10500 12500 10580 12520
rect 10500 12140 10520 12500
rect 10560 12140 10580 12500
rect 10500 12120 10580 12140
rect 10610 12120 10730 12520
rect 10760 12500 10840 12520
rect 10760 12140 10780 12500
rect 10820 12140 10840 12500
rect 10760 12120 10840 12140
rect 10870 12120 10940 12520
rect 11000 12300 11070 12320
rect 11000 12140 11010 12300
rect 11050 12140 11070 12300
rect 11000 12120 11070 12140
rect 11100 12300 11180 12320
rect 11100 12140 11120 12300
rect 11160 12140 11180 12300
rect 11100 12120 11180 12140
rect 11210 12300 11280 12320
rect 11210 12140 11230 12300
rect 11270 12140 11280 12300
rect 11210 12120 11280 12140
rect 11390 12120 11460 12520
rect 11490 12500 11570 12520
rect 11490 12140 11510 12500
rect 11550 12140 11570 12500
rect 11490 12120 11570 12140
rect 11600 12120 11720 12520
rect 11750 12500 11830 12520
rect 11750 12140 11770 12500
rect 11810 12140 11830 12500
rect 11750 12120 11830 12140
rect 11860 12120 11930 12520
rect 11990 12300 12060 12320
rect 11990 12140 12000 12300
rect 12040 12140 12060 12300
rect 11990 12120 12060 12140
rect 12090 12300 12170 12320
rect 12090 12140 12110 12300
rect 12150 12140 12170 12300
rect 12090 12120 12170 12140
rect 12200 12300 12270 12320
rect 12200 12140 12220 12300
rect 12260 12140 12270 12300
rect 12200 12120 12270 12140
rect 12390 12120 12460 12520
rect 12490 12500 12570 12520
rect 12490 12140 12510 12500
rect 12550 12140 12570 12500
rect 12490 12120 12570 12140
rect 12600 12120 12720 12520
rect 12750 12500 12830 12520
rect 12750 12140 12770 12500
rect 12810 12140 12830 12500
rect 12750 12120 12830 12140
rect 12860 12120 12930 12520
rect 13340 12580 13410 12600
rect 13340 12420 13350 12580
rect 13390 12420 13410 12580
rect 13340 12400 13410 12420
rect 13440 12580 13510 12600
rect 13440 12420 13460 12580
rect 13500 12420 13510 12580
rect 13440 12400 13510 12420
rect 13570 12580 13640 12600
rect 13570 12420 13580 12580
rect 13620 12420 13640 12580
rect 13570 12400 13640 12420
rect 13670 12580 13750 12600
rect 13670 12420 13690 12580
rect 13730 12420 13750 12580
rect 13670 12400 13750 12420
rect 13780 12580 13850 12600
rect 13780 12420 13800 12580
rect 13840 12420 13850 12580
rect 13780 12400 13850 12420
rect 13910 12580 13980 12600
rect 13910 12420 13920 12580
rect 13960 12420 13980 12580
rect 13910 12400 13980 12420
rect 14010 12580 14090 12600
rect 14010 12420 14030 12580
rect 14070 12420 14090 12580
rect 14010 12400 14090 12420
rect 14120 12580 14200 12600
rect 14120 12420 14140 12580
rect 14180 12420 14200 12580
rect 14120 12400 14200 12420
rect 14230 12580 14310 12600
rect 14230 12420 14250 12580
rect 14290 12420 14310 12580
rect 14230 12400 14310 12420
rect 14340 12580 14410 12600
rect 14340 12420 14360 12580
rect 14400 12420 14410 12580
rect 14340 12400 14410 12420
rect 14470 12580 14540 12600
rect 14470 12420 14480 12580
rect 14520 12420 14540 12580
rect 14470 12400 14540 12420
rect 14570 12580 14650 12600
rect 14570 12420 14590 12580
rect 14630 12420 14650 12580
rect 14570 12400 14650 12420
rect 14680 12580 14760 12600
rect 14680 12420 14700 12580
rect 14740 12420 14760 12580
rect 14680 12400 14760 12420
rect 14790 12580 14870 12600
rect 14790 12420 14810 12580
rect 14850 12420 14870 12580
rect 14790 12400 14870 12420
rect 14900 12580 14980 12600
rect 14900 12420 14920 12580
rect 14960 12420 14980 12580
rect 14900 12400 14980 12420
rect 15010 12580 15090 12600
rect 15010 12420 15030 12580
rect 15070 12420 15090 12580
rect 15010 12400 15090 12420
rect 15120 12580 15200 12600
rect 15120 12420 15140 12580
rect 15180 12420 15200 12580
rect 15120 12400 15200 12420
rect 15230 12580 15310 12600
rect 15230 12420 15250 12580
rect 15290 12420 15310 12580
rect 15230 12400 15310 12420
rect 15340 12580 15410 12600
rect 15340 12420 15360 12580
rect 15400 12420 15410 12580
rect 15340 12400 15410 12420
rect 15530 12580 15600 12600
rect 15530 12420 15540 12580
rect 15580 12420 15600 12580
rect 15530 12400 15600 12420
rect 15630 12580 15710 12600
rect 15630 12420 15650 12580
rect 15690 12420 15710 12580
rect 15630 12400 15710 12420
rect 15740 12580 15820 12600
rect 15740 12420 15760 12580
rect 15800 12420 15820 12580
rect 15740 12400 15820 12420
rect 15850 12580 15930 12600
rect 15850 12420 15870 12580
rect 15910 12420 15930 12580
rect 15850 12400 15930 12420
rect 15960 12580 16040 12600
rect 15960 12420 15980 12580
rect 16020 12420 16040 12580
rect 15960 12400 16040 12420
rect 16070 12580 16150 12600
rect 16070 12420 16090 12580
rect 16130 12420 16150 12580
rect 16070 12400 16150 12420
rect 16180 12580 16260 12600
rect 16180 12420 16200 12580
rect 16240 12420 16260 12580
rect 16180 12400 16260 12420
rect 16290 12580 16370 12600
rect 16290 12420 16310 12580
rect 16350 12420 16370 12580
rect 16290 12400 16370 12420
rect 16400 12580 16480 12600
rect 16400 12420 16420 12580
rect 16460 12420 16480 12580
rect 16400 12400 16480 12420
rect 16510 12580 16590 12600
rect 16510 12420 16530 12580
rect 16570 12420 16590 12580
rect 16510 12400 16590 12420
rect 16620 12580 16700 12600
rect 16620 12420 16640 12580
rect 16680 12420 16700 12580
rect 16620 12400 16700 12420
rect 16730 12580 16810 12600
rect 16730 12420 16750 12580
rect 16790 12420 16810 12580
rect 16730 12400 16810 12420
rect 16840 12580 16920 12600
rect 16840 12420 16860 12580
rect 16900 12420 16920 12580
rect 16840 12400 16920 12420
rect 16950 12580 17030 12600
rect 16950 12420 16970 12580
rect 17010 12420 17030 12580
rect 16950 12400 17030 12420
rect 17060 12580 17140 12600
rect 17060 12420 17080 12580
rect 17120 12420 17140 12580
rect 17060 12400 17140 12420
rect 17170 12580 17250 12600
rect 17170 12420 17190 12580
rect 17230 12420 17250 12580
rect 17170 12400 17250 12420
rect 17280 12580 17350 12600
rect 17280 12420 17300 12580
rect 17340 12420 17350 12580
rect 17280 12400 17350 12420
rect 17480 12580 17550 12600
rect 17480 12420 17490 12580
rect 17530 12420 17550 12580
rect 17480 12400 17550 12420
rect 17580 12580 17660 12600
rect 17580 12420 17600 12580
rect 17640 12420 17660 12580
rect 17580 12400 17660 12420
rect 17690 12580 17770 12600
rect 17690 12420 17710 12580
rect 17750 12420 17770 12580
rect 17690 12400 17770 12420
rect 17800 12580 17880 12600
rect 17800 12420 17820 12580
rect 17860 12420 17880 12580
rect 17800 12400 17880 12420
rect 17910 12580 17990 12600
rect 17910 12420 17930 12580
rect 17970 12420 17990 12580
rect 17910 12400 17990 12420
rect 18020 12580 18100 12600
rect 18020 12420 18040 12580
rect 18080 12420 18100 12580
rect 18020 12400 18100 12420
rect 18130 12580 18210 12600
rect 18130 12420 18150 12580
rect 18190 12420 18210 12580
rect 18130 12400 18210 12420
rect 18240 12580 18320 12600
rect 18240 12420 18260 12580
rect 18300 12420 18320 12580
rect 18240 12400 18320 12420
rect 18350 12580 18430 12600
rect 18350 12420 18370 12580
rect 18410 12420 18430 12580
rect 18350 12400 18430 12420
rect 18460 12580 18540 12600
rect 18460 12420 18480 12580
rect 18520 12420 18540 12580
rect 18460 12400 18540 12420
rect 18570 12580 18650 12600
rect 18570 12420 18590 12580
rect 18630 12420 18650 12580
rect 18570 12400 18650 12420
rect 18680 12580 18760 12600
rect 18680 12420 18700 12580
rect 18740 12420 18760 12580
rect 18680 12400 18760 12420
rect 18790 12580 18870 12600
rect 18790 12420 18810 12580
rect 18850 12420 18870 12580
rect 18790 12400 18870 12420
rect 18900 12580 18980 12600
rect 18900 12420 18920 12580
rect 18960 12420 18980 12580
rect 18900 12400 18980 12420
rect 19010 12580 19090 12600
rect 19010 12420 19030 12580
rect 19070 12420 19090 12580
rect 19010 12400 19090 12420
rect 19120 12580 19200 12600
rect 19120 12420 19140 12580
rect 19180 12420 19200 12580
rect 19120 12400 19200 12420
rect 19230 12580 19310 12600
rect 19230 12420 19250 12580
rect 19290 12420 19310 12580
rect 19230 12400 19310 12420
rect 19340 12580 19420 12600
rect 19340 12420 19360 12580
rect 19400 12420 19420 12580
rect 19340 12400 19420 12420
rect 19450 12580 19530 12600
rect 19450 12420 19470 12580
rect 19510 12420 19530 12580
rect 19450 12400 19530 12420
rect 19560 12580 19640 12600
rect 19560 12420 19580 12580
rect 19620 12420 19640 12580
rect 19560 12400 19640 12420
rect 19670 12580 19750 12600
rect 19670 12420 19690 12580
rect 19730 12420 19750 12580
rect 19670 12400 19750 12420
rect 19780 12580 19860 12600
rect 19780 12420 19800 12580
rect 19840 12420 19860 12580
rect 19780 12400 19860 12420
rect 19890 12580 19970 12600
rect 19890 12420 19910 12580
rect 19950 12420 19970 12580
rect 19890 12400 19970 12420
rect 20000 12580 20080 12600
rect 20000 12420 20020 12580
rect 20060 12420 20080 12580
rect 20000 12400 20080 12420
rect 20110 12580 20190 12600
rect 20110 12420 20130 12580
rect 20170 12420 20190 12580
rect 20110 12400 20190 12420
rect 20220 12580 20300 12600
rect 20220 12420 20240 12580
rect 20280 12420 20300 12580
rect 20220 12400 20300 12420
rect 20330 12580 20410 12600
rect 20330 12420 20350 12580
rect 20390 12420 20410 12580
rect 20330 12400 20410 12420
rect 20440 12580 20520 12600
rect 20440 12420 20460 12580
rect 20500 12420 20520 12580
rect 20440 12400 20520 12420
rect 20550 12580 20630 12600
rect 20550 12420 20570 12580
rect 20610 12420 20630 12580
rect 20550 12400 20630 12420
rect 20660 12580 20740 12600
rect 20660 12420 20680 12580
rect 20720 12420 20740 12580
rect 20660 12400 20740 12420
rect 20770 12580 20850 12600
rect 20770 12420 20790 12580
rect 20830 12420 20850 12580
rect 20770 12400 20850 12420
rect 20880 12580 20960 12600
rect 20880 12420 20900 12580
rect 20940 12420 20960 12580
rect 20880 12400 20960 12420
rect 20990 12580 21060 12600
rect 20990 12420 21010 12580
rect 21050 12420 21060 12580
rect 20990 12400 21060 12420
rect 12990 12300 13060 12320
rect 12990 12140 13000 12300
rect 13040 12140 13060 12300
rect 12990 12120 13060 12140
rect 13090 12300 13170 12320
rect 13090 12140 13110 12300
rect 13150 12140 13170 12300
rect 13090 12120 13170 12140
rect 13200 12300 13270 12320
rect 13200 12140 13220 12300
rect 13260 12140 13270 12300
rect 13200 12120 13270 12140
rect 8800 12080 8870 12100
rect 7850 11280 7920 11300
rect 7850 11120 7860 11280
rect 7900 11120 7920 11280
rect 7850 11100 7920 11120
rect 7950 11280 8030 11300
rect 7950 11120 7970 11280
rect 8010 11120 8030 11280
rect 7950 11100 8030 11120
rect 8060 11280 8180 11300
rect 8060 11120 8100 11280
rect 8140 11120 8180 11280
rect 8060 11100 8180 11120
rect 8210 11280 8290 11300
rect 8210 11120 8230 11280
rect 8270 11120 8290 11280
rect 8210 11100 8290 11120
rect 8320 11280 8390 11300
rect 8320 11120 8340 11280
rect 8380 11120 8390 11280
rect 8320 11100 8390 11120
rect 7280 10910 7350 10930
rect 7280 10750 7290 10910
rect 7330 10750 7350 10910
rect 7280 10730 7350 10750
rect 7380 10910 7460 10930
rect 7380 10750 7400 10910
rect 7440 10750 7460 10910
rect 7380 10730 7460 10750
rect 7490 10910 7560 10930
rect 7490 10750 7510 10910
rect 7550 10750 7560 10910
rect 7490 10730 7560 10750
rect 8640 10960 8710 10980
rect 8640 10600 8650 10960
rect 8690 10600 8710 10960
rect 8640 10580 8710 10600
rect 8740 10960 8860 10980
rect 8740 10600 8780 10960
rect 8820 10600 8860 10960
rect 8740 10580 8860 10600
rect 8890 10960 8960 10980
rect 8890 10600 8910 10960
rect 8950 10600 8960 10960
rect 9860 10910 9930 10930
rect 9860 10750 9870 10910
rect 9910 10750 9930 10910
rect 9860 10730 9930 10750
rect 9960 10910 10040 10930
rect 9960 10750 9980 10910
rect 10020 10750 10040 10910
rect 9960 10730 10040 10750
rect 10070 10910 10140 10930
rect 10070 10750 10090 10910
rect 10130 10750 10140 10910
rect 10070 10730 10140 10750
rect 8890 10580 8960 10600
rect 9020 10650 9090 10670
rect 9020 10490 9030 10650
rect 9070 10490 9090 10650
rect 9020 10470 9090 10490
rect 9120 10650 9190 10670
rect 9120 10490 9140 10650
rect 9180 10490 9190 10650
rect 9120 10470 9190 10490
rect 9280 10650 9350 10670
rect 9280 10490 9290 10650
rect 9330 10490 9350 10650
rect 9280 10470 9350 10490
rect 9380 10650 9450 10670
rect 9380 10490 9400 10650
rect 9440 10490 9450 10650
rect 9380 10470 9450 10490
rect 9530 10650 9600 10670
rect 9530 10490 9540 10650
rect 9580 10490 9600 10650
rect 9530 10470 9600 10490
rect 9630 10650 9700 10670
rect 9630 10490 9650 10650
rect 9690 10490 9700 10650
rect 9630 10470 9700 10490
rect 10400 10530 10470 10930
rect 10500 10910 10580 10930
rect 10500 10550 10520 10910
rect 10560 10550 10580 10910
rect 10500 10530 10580 10550
rect 10610 10530 10730 10930
rect 10760 10910 10840 10930
rect 10760 10550 10780 10910
rect 10820 10550 10840 10910
rect 10760 10530 10840 10550
rect 10870 10530 10940 10930
rect 11000 10910 11070 10930
rect 11000 10750 11010 10910
rect 11050 10750 11070 10910
rect 11000 10730 11070 10750
rect 11100 10910 11180 10930
rect 11100 10750 11120 10910
rect 11160 10750 11180 10910
rect 11100 10730 11180 10750
rect 11210 10910 11280 10930
rect 11210 10750 11230 10910
rect 11270 10750 11280 10910
rect 11210 10730 11280 10750
rect 11390 10530 11460 10930
rect 11490 10910 11570 10930
rect 11490 10550 11510 10910
rect 11550 10550 11570 10910
rect 11490 10530 11570 10550
rect 11600 10530 11720 10930
rect 11750 10910 11830 10930
rect 11750 10550 11770 10910
rect 11810 10550 11830 10910
rect 11750 10530 11830 10550
rect 11860 10530 11930 10930
rect 11990 10910 12060 10930
rect 11990 10750 12000 10910
rect 12040 10750 12060 10910
rect 11990 10730 12060 10750
rect 12090 10910 12170 10930
rect 12090 10750 12110 10910
rect 12150 10750 12170 10910
rect 12090 10730 12170 10750
rect 12200 10910 12270 10930
rect 12200 10750 12220 10910
rect 12260 10750 12270 10910
rect 12200 10730 12270 10750
rect 12390 10530 12460 10930
rect 12490 10910 12570 10930
rect 12490 10550 12510 10910
rect 12550 10550 12570 10910
rect 12490 10530 12570 10550
rect 12600 10530 12720 10930
rect 12750 10910 12830 10930
rect 12750 10550 12770 10910
rect 12810 10550 12830 10910
rect 12750 10530 12830 10550
rect 12860 10530 12930 10930
rect 12990 10910 13060 10930
rect 12990 10750 13000 10910
rect 13040 10750 13060 10910
rect 12990 10730 13060 10750
rect 13090 10910 13170 10930
rect 13090 10750 13110 10910
rect 13150 10750 13170 10910
rect 13090 10730 13170 10750
rect 13200 10910 13270 10930
rect 13200 10750 13220 10910
rect 13260 10750 13270 10910
rect 13200 10730 13270 10750
rect 13330 10630 13400 10650
rect 13330 10470 13340 10630
rect 13380 10470 13400 10630
rect 13330 10450 13400 10470
rect 13430 10630 13500 10650
rect 13430 10470 13450 10630
rect 13490 10470 13500 10630
rect 13430 10450 13500 10470
rect 13560 10630 13630 10650
rect 13560 10470 13570 10630
rect 13610 10470 13630 10630
rect 13560 10450 13630 10470
rect 13660 10630 13740 10650
rect 13660 10470 13680 10630
rect 13720 10470 13740 10630
rect 13660 10450 13740 10470
rect 13770 10630 13840 10650
rect 13770 10470 13790 10630
rect 13830 10470 13840 10630
rect 13770 10450 13840 10470
rect 13900 10630 13970 10650
rect 13900 10470 13910 10630
rect 13950 10470 13970 10630
rect 13900 10450 13970 10470
rect 14000 10630 14080 10650
rect 14000 10470 14020 10630
rect 14060 10470 14080 10630
rect 14000 10450 14080 10470
rect 14110 10630 14190 10650
rect 14110 10470 14130 10630
rect 14170 10470 14190 10630
rect 14110 10450 14190 10470
rect 14220 10630 14300 10650
rect 14220 10470 14240 10630
rect 14280 10470 14300 10630
rect 14220 10450 14300 10470
rect 14330 10630 14400 10650
rect 14330 10470 14350 10630
rect 14390 10470 14400 10630
rect 14330 10450 14400 10470
rect 14460 10630 14530 10650
rect 14460 10470 14470 10630
rect 14510 10470 14530 10630
rect 14460 10450 14530 10470
rect 14560 10630 14640 10650
rect 14560 10470 14580 10630
rect 14620 10470 14640 10630
rect 14560 10450 14640 10470
rect 14670 10630 14750 10650
rect 14670 10470 14690 10630
rect 14730 10470 14750 10630
rect 14670 10450 14750 10470
rect 14780 10630 14860 10650
rect 14780 10470 14800 10630
rect 14840 10470 14860 10630
rect 14780 10450 14860 10470
rect 14890 10630 14970 10650
rect 14890 10470 14910 10630
rect 14950 10470 14970 10630
rect 14890 10450 14970 10470
rect 15000 10630 15080 10650
rect 15000 10470 15020 10630
rect 15060 10470 15080 10630
rect 15000 10450 15080 10470
rect 15110 10630 15190 10650
rect 15110 10470 15130 10630
rect 15170 10470 15190 10630
rect 15110 10450 15190 10470
rect 15220 10630 15300 10650
rect 15220 10470 15240 10630
rect 15280 10470 15300 10630
rect 15220 10450 15300 10470
rect 15330 10630 15400 10650
rect 15330 10470 15350 10630
rect 15390 10470 15400 10630
rect 15330 10450 15400 10470
rect 15520 10630 15590 10650
rect 15520 10470 15530 10630
rect 15570 10470 15590 10630
rect 15520 10450 15590 10470
rect 15620 10630 15700 10650
rect 15620 10470 15640 10630
rect 15680 10470 15700 10630
rect 15620 10450 15700 10470
rect 15730 10630 15810 10650
rect 15730 10470 15750 10630
rect 15790 10470 15810 10630
rect 15730 10450 15810 10470
rect 15840 10630 15920 10650
rect 15840 10470 15860 10630
rect 15900 10470 15920 10630
rect 15840 10450 15920 10470
rect 15950 10630 16030 10650
rect 15950 10470 15970 10630
rect 16010 10470 16030 10630
rect 15950 10450 16030 10470
rect 16060 10630 16140 10650
rect 16060 10470 16080 10630
rect 16120 10470 16140 10630
rect 16060 10450 16140 10470
rect 16170 10630 16250 10650
rect 16170 10470 16190 10630
rect 16230 10470 16250 10630
rect 16170 10450 16250 10470
rect 16280 10630 16360 10650
rect 16280 10470 16300 10630
rect 16340 10470 16360 10630
rect 16280 10450 16360 10470
rect 16390 10630 16470 10650
rect 16390 10470 16410 10630
rect 16450 10470 16470 10630
rect 16390 10450 16470 10470
rect 16500 10630 16580 10650
rect 16500 10470 16520 10630
rect 16560 10470 16580 10630
rect 16500 10450 16580 10470
rect 16610 10630 16690 10650
rect 16610 10470 16630 10630
rect 16670 10470 16690 10630
rect 16610 10450 16690 10470
rect 16720 10630 16800 10650
rect 16720 10470 16740 10630
rect 16780 10470 16800 10630
rect 16720 10450 16800 10470
rect 16830 10630 16910 10650
rect 16830 10470 16850 10630
rect 16890 10470 16910 10630
rect 16830 10450 16910 10470
rect 16940 10630 17020 10650
rect 16940 10470 16960 10630
rect 17000 10470 17020 10630
rect 16940 10450 17020 10470
rect 17050 10630 17130 10650
rect 17050 10470 17070 10630
rect 17110 10470 17130 10630
rect 17050 10450 17130 10470
rect 17160 10630 17240 10650
rect 17160 10470 17180 10630
rect 17220 10470 17240 10630
rect 17160 10450 17240 10470
rect 17270 10630 17340 10650
rect 17270 10470 17290 10630
rect 17330 10470 17340 10630
rect 17270 10450 17340 10470
rect 17470 10630 17540 10650
rect 17470 10470 17480 10630
rect 17520 10470 17540 10630
rect 17470 10450 17540 10470
rect 17570 10630 17650 10650
rect 17570 10470 17590 10630
rect 17630 10470 17650 10630
rect 17570 10450 17650 10470
rect 17680 10630 17760 10650
rect 17680 10470 17700 10630
rect 17740 10470 17760 10630
rect 17680 10450 17760 10470
rect 17790 10630 17870 10650
rect 17790 10470 17810 10630
rect 17850 10470 17870 10630
rect 17790 10450 17870 10470
rect 17900 10630 17980 10650
rect 17900 10470 17920 10630
rect 17960 10470 17980 10630
rect 17900 10450 17980 10470
rect 18010 10630 18090 10650
rect 18010 10470 18030 10630
rect 18070 10470 18090 10630
rect 18010 10450 18090 10470
rect 18120 10630 18200 10650
rect 18120 10470 18140 10630
rect 18180 10470 18200 10630
rect 18120 10450 18200 10470
rect 18230 10630 18310 10650
rect 18230 10470 18250 10630
rect 18290 10470 18310 10630
rect 18230 10450 18310 10470
rect 18340 10630 18420 10650
rect 18340 10470 18360 10630
rect 18400 10470 18420 10630
rect 18340 10450 18420 10470
rect 18450 10630 18530 10650
rect 18450 10470 18470 10630
rect 18510 10470 18530 10630
rect 18450 10450 18530 10470
rect 18560 10630 18640 10650
rect 18560 10470 18580 10630
rect 18620 10470 18640 10630
rect 18560 10450 18640 10470
rect 18670 10630 18750 10650
rect 18670 10470 18690 10630
rect 18730 10470 18750 10630
rect 18670 10450 18750 10470
rect 18780 10630 18860 10650
rect 18780 10470 18800 10630
rect 18840 10470 18860 10630
rect 18780 10450 18860 10470
rect 18890 10630 18970 10650
rect 18890 10470 18910 10630
rect 18950 10470 18970 10630
rect 18890 10450 18970 10470
rect 19000 10630 19080 10650
rect 19000 10470 19020 10630
rect 19060 10470 19080 10630
rect 19000 10450 19080 10470
rect 19110 10630 19190 10650
rect 19110 10470 19130 10630
rect 19170 10470 19190 10630
rect 19110 10450 19190 10470
rect 19220 10630 19300 10650
rect 19220 10470 19240 10630
rect 19280 10470 19300 10630
rect 19220 10450 19300 10470
rect 19330 10630 19410 10650
rect 19330 10470 19350 10630
rect 19390 10470 19410 10630
rect 19330 10450 19410 10470
rect 19440 10630 19520 10650
rect 19440 10470 19460 10630
rect 19500 10470 19520 10630
rect 19440 10450 19520 10470
rect 19550 10630 19630 10650
rect 19550 10470 19570 10630
rect 19610 10470 19630 10630
rect 19550 10450 19630 10470
rect 19660 10630 19740 10650
rect 19660 10470 19680 10630
rect 19720 10470 19740 10630
rect 19660 10450 19740 10470
rect 19770 10630 19850 10650
rect 19770 10470 19790 10630
rect 19830 10470 19850 10630
rect 19770 10450 19850 10470
rect 19880 10630 19960 10650
rect 19880 10470 19900 10630
rect 19940 10470 19960 10630
rect 19880 10450 19960 10470
rect 19990 10630 20070 10650
rect 19990 10470 20010 10630
rect 20050 10470 20070 10630
rect 19990 10450 20070 10470
rect 20100 10630 20180 10650
rect 20100 10470 20120 10630
rect 20160 10470 20180 10630
rect 20100 10450 20180 10470
rect 20210 10630 20290 10650
rect 20210 10470 20230 10630
rect 20270 10470 20290 10630
rect 20210 10450 20290 10470
rect 20320 10630 20400 10650
rect 20320 10470 20340 10630
rect 20380 10470 20400 10630
rect 20320 10450 20400 10470
rect 20430 10630 20510 10650
rect 20430 10470 20450 10630
rect 20490 10470 20510 10630
rect 20430 10450 20510 10470
rect 20540 10630 20620 10650
rect 20540 10470 20560 10630
rect 20600 10470 20620 10630
rect 20540 10450 20620 10470
rect 20650 10630 20730 10650
rect 20650 10470 20670 10630
rect 20710 10470 20730 10630
rect 20650 10450 20730 10470
rect 20760 10630 20840 10650
rect 20760 10470 20780 10630
rect 20820 10470 20840 10630
rect 20760 10450 20840 10470
rect 20870 10630 20950 10650
rect 20870 10470 20890 10630
rect 20930 10470 20950 10630
rect 20870 10450 20950 10470
rect 20980 10630 21050 10650
rect 20980 10470 21000 10630
rect 21040 10470 21050 10630
rect 20980 10450 21050 10470
rect 13630 4120 13700 4140
rect 9870 3790 9940 3810
rect 9870 3230 9880 3790
rect 9920 3230 9940 3790
rect 9870 3210 9940 3230
rect 9970 3790 10050 3810
rect 9970 3230 9990 3790
rect 10030 3230 10050 3790
rect 9970 3210 10050 3230
rect 10080 3790 10160 3810
rect 10080 3230 10100 3790
rect 10140 3230 10160 3790
rect 10080 3210 10160 3230
rect 10190 3790 10270 3810
rect 10190 3230 10210 3790
rect 10250 3230 10270 3790
rect 10190 3210 10270 3230
rect 10300 3790 10380 3810
rect 10300 3230 10320 3790
rect 10360 3230 10380 3790
rect 10300 3210 10380 3230
rect 10410 3790 10490 3810
rect 10410 3230 10430 3790
rect 10470 3230 10490 3790
rect 10410 3210 10490 3230
rect 10520 3790 10600 3810
rect 10520 3230 10540 3790
rect 10580 3230 10600 3790
rect 10520 3210 10600 3230
rect 10630 3790 10710 3810
rect 10630 3230 10650 3790
rect 10690 3230 10710 3790
rect 10630 3210 10710 3230
rect 10740 3790 10820 3810
rect 10740 3230 10760 3790
rect 10800 3230 10820 3790
rect 10740 3210 10820 3230
rect 10850 3790 10930 3810
rect 10850 3230 10870 3790
rect 10910 3230 10930 3790
rect 10850 3210 10930 3230
rect 10960 3790 11040 3810
rect 10960 3230 10980 3790
rect 11020 3230 11040 3790
rect 10960 3210 11040 3230
rect 11070 3790 11150 3810
rect 11070 3230 11090 3790
rect 11130 3230 11150 3790
rect 11070 3210 11150 3230
rect 11180 3790 11260 3810
rect 11180 3230 11200 3790
rect 11240 3230 11260 3790
rect 11180 3210 11260 3230
rect 11290 3790 11370 3810
rect 11290 3230 11310 3790
rect 11350 3230 11370 3790
rect 11290 3210 11370 3230
rect 11400 3790 11480 3810
rect 11400 3230 11420 3790
rect 11460 3230 11480 3790
rect 11400 3210 11480 3230
rect 11510 3790 11590 3810
rect 11510 3230 11530 3790
rect 11570 3230 11590 3790
rect 11510 3210 11590 3230
rect 11620 3790 11700 3810
rect 11620 3230 11640 3790
rect 11680 3230 11700 3790
rect 11620 3210 11700 3230
rect 11730 3790 11810 3810
rect 11730 3230 11750 3790
rect 11790 3230 11810 3790
rect 11730 3210 11810 3230
rect 11840 3790 11920 3810
rect 11840 3230 11860 3790
rect 11900 3230 11920 3790
rect 11840 3210 11920 3230
rect 11950 3790 12030 3810
rect 11950 3230 11970 3790
rect 12010 3230 12030 3790
rect 11950 3210 12030 3230
rect 12060 3790 12140 3810
rect 12060 3230 12080 3790
rect 12120 3230 12140 3790
rect 12060 3210 12140 3230
rect 12170 3790 12250 3810
rect 12170 3230 12190 3790
rect 12230 3230 12250 3790
rect 12170 3210 12250 3230
rect 12280 3790 12360 3810
rect 12280 3230 12300 3790
rect 12340 3230 12360 3790
rect 12280 3210 12360 3230
rect 12390 3790 12470 3810
rect 12390 3230 12410 3790
rect 12450 3230 12470 3790
rect 12390 3210 12470 3230
rect 12500 3790 12580 3810
rect 12500 3230 12520 3790
rect 12560 3230 12580 3790
rect 12500 3210 12580 3230
rect 12610 3790 12690 3810
rect 12610 3230 12630 3790
rect 12670 3230 12690 3790
rect 12610 3210 12690 3230
rect 12720 3790 12800 3810
rect 12720 3230 12740 3790
rect 12780 3230 12800 3790
rect 12720 3210 12800 3230
rect 12830 3790 12910 3810
rect 12830 3230 12850 3790
rect 12890 3230 12910 3790
rect 12830 3210 12910 3230
rect 12940 3790 13020 3810
rect 12940 3230 12960 3790
rect 13000 3230 13020 3790
rect 12940 3210 13020 3230
rect 13050 3790 13130 3810
rect 13050 3230 13070 3790
rect 13110 3230 13130 3790
rect 13050 3210 13130 3230
rect 13160 3790 13230 3810
rect 13160 3230 13180 3790
rect 13220 3230 13230 3790
rect 13630 3560 13640 4120
rect 13680 3560 13700 4120
rect 13630 3540 13700 3560
rect 13730 4120 13810 4140
rect 13730 3560 13750 4120
rect 13790 3560 13810 4120
rect 13730 3540 13810 3560
rect 13840 4120 13920 4140
rect 13840 3560 13860 4120
rect 13900 3560 13920 4120
rect 13840 3540 13920 3560
rect 13950 4120 14030 4140
rect 13950 3560 13970 4120
rect 14010 3560 14030 4120
rect 13950 3540 14030 3560
rect 14060 4120 14140 4140
rect 14060 3560 14080 4120
rect 14120 3560 14140 4120
rect 14060 3540 14140 3560
rect 14170 4120 14250 4140
rect 14170 3560 14190 4120
rect 14230 3560 14250 4120
rect 14170 3540 14250 3560
rect 14280 4120 14360 4140
rect 14280 3560 14300 4120
rect 14340 3560 14360 4120
rect 14280 3540 14360 3560
rect 14390 4120 14470 4140
rect 14390 3560 14410 4120
rect 14450 3560 14470 4120
rect 14390 3540 14470 3560
rect 14500 4120 14580 4140
rect 14500 3560 14520 4120
rect 14560 3560 14580 4120
rect 14500 3540 14580 3560
rect 14610 4120 14690 4140
rect 14610 3560 14630 4120
rect 14670 3560 14690 4120
rect 14610 3540 14690 3560
rect 14720 4120 14800 4140
rect 14720 3560 14740 4120
rect 14780 3560 14800 4120
rect 14720 3540 14800 3560
rect 14830 4120 14910 4140
rect 14830 3560 14850 4120
rect 14890 3560 14910 4120
rect 14830 3540 14910 3560
rect 14940 4120 15020 4140
rect 14940 3560 14960 4120
rect 15000 3560 15020 4120
rect 14940 3540 15020 3560
rect 15050 4120 15130 4140
rect 15050 3560 15070 4120
rect 15110 3560 15130 4120
rect 15050 3540 15130 3560
rect 15160 4120 15240 4140
rect 15160 3560 15180 4120
rect 15220 3560 15240 4120
rect 15160 3540 15240 3560
rect 15270 4120 15350 4140
rect 15270 3560 15290 4120
rect 15330 3560 15350 4120
rect 15270 3540 15350 3560
rect 15380 4120 15460 4140
rect 15380 3560 15400 4120
rect 15440 3560 15460 4120
rect 15380 3540 15460 3560
rect 15490 4120 15570 4140
rect 15490 3560 15510 4120
rect 15550 3560 15570 4120
rect 15490 3540 15570 3560
rect 15600 4120 15680 4140
rect 15600 3560 15620 4120
rect 15660 3560 15680 4120
rect 15600 3540 15680 3560
rect 15710 4120 15790 4140
rect 15710 3560 15730 4120
rect 15770 3560 15790 4120
rect 15710 3540 15790 3560
rect 15820 4120 15900 4140
rect 15820 3560 15840 4120
rect 15880 3560 15900 4120
rect 15820 3540 15900 3560
rect 15930 4120 16010 4140
rect 15930 3560 15950 4120
rect 15990 3560 16010 4120
rect 15930 3540 16010 3560
rect 16040 4120 16120 4140
rect 16040 3560 16060 4120
rect 16100 3560 16120 4120
rect 16040 3540 16120 3560
rect 16150 4120 16230 4140
rect 16150 3560 16170 4120
rect 16210 3560 16230 4120
rect 16150 3540 16230 3560
rect 16260 4120 16340 4140
rect 16260 3560 16280 4120
rect 16320 3560 16340 4120
rect 16260 3540 16340 3560
rect 16370 4120 16450 4140
rect 16370 3560 16390 4120
rect 16430 3560 16450 4120
rect 16370 3540 16450 3560
rect 16480 4120 16560 4140
rect 16480 3560 16500 4120
rect 16540 3560 16560 4120
rect 16480 3540 16560 3560
rect 16590 4120 16670 4140
rect 16590 3560 16610 4120
rect 16650 3560 16670 4120
rect 16590 3540 16670 3560
rect 16700 4120 16780 4140
rect 16700 3560 16720 4120
rect 16760 3560 16780 4120
rect 16700 3540 16780 3560
rect 16810 4120 16890 4140
rect 16810 3560 16830 4120
rect 16870 3560 16890 4120
rect 16810 3540 16890 3560
rect 16920 4120 16990 4140
rect 16920 3560 16940 4120
rect 16980 3560 16990 4120
rect 16920 3540 16990 3560
rect 13160 3210 13230 3230
rect 24350 2760 25350 2770
rect 24350 2720 24370 2760
rect 25330 2720 25350 2760
rect 24350 2700 25350 2720
rect 24350 2650 25350 2670
rect 24350 2610 24370 2650
rect 25330 2610 25350 2650
rect 24350 2590 25350 2610
rect 24350 2540 25350 2560
rect 24350 2500 24370 2540
rect 25330 2500 25350 2540
rect 24350 2480 25350 2500
rect 24350 2430 25350 2450
rect 24350 2390 24370 2430
rect 25330 2390 25350 2430
rect 24350 2370 25350 2390
rect 24350 2320 25350 2340
rect 24350 2280 24370 2320
rect 25330 2280 25350 2320
rect 24350 2260 25350 2280
rect 24350 2210 25350 2230
rect 24350 2170 24370 2210
rect 25330 2170 25350 2210
rect 24350 2150 25350 2170
rect 24350 2100 25350 2120
rect 24350 2060 24370 2100
rect 25330 2060 25350 2100
rect 24350 2050 25350 2060
rect 9890 1310 9960 1330
rect 9890 750 9900 1310
rect 9940 750 9960 1310
rect 9890 730 9960 750
rect 9990 1310 10070 1330
rect 9990 750 10010 1310
rect 10050 750 10070 1310
rect 9990 730 10070 750
rect 10100 1310 10180 1330
rect 10100 750 10120 1310
rect 10160 750 10180 1310
rect 10100 730 10180 750
rect 10210 1310 10290 1330
rect 10210 750 10230 1310
rect 10270 750 10290 1310
rect 10210 730 10290 750
rect 10320 1310 10400 1330
rect 10320 750 10340 1310
rect 10380 750 10400 1310
rect 10320 730 10400 750
rect 10430 1310 10510 1330
rect 10430 750 10450 1310
rect 10490 750 10510 1310
rect 10430 730 10510 750
rect 10540 1310 10620 1330
rect 10540 750 10560 1310
rect 10600 750 10620 1310
rect 10540 730 10620 750
rect 10650 1310 10730 1330
rect 10650 750 10670 1310
rect 10710 750 10730 1310
rect 10650 730 10730 750
rect 10760 1310 10840 1330
rect 10760 750 10780 1310
rect 10820 750 10840 1310
rect 10760 730 10840 750
rect 10870 1310 10950 1330
rect 10870 750 10890 1310
rect 10930 750 10950 1310
rect 10870 730 10950 750
rect 10980 1310 11060 1330
rect 10980 750 11000 1310
rect 11040 750 11060 1310
rect 10980 730 11060 750
rect 11090 1310 11170 1330
rect 11090 750 11110 1310
rect 11150 750 11170 1310
rect 11090 730 11170 750
rect 11200 1310 11280 1330
rect 11200 750 11220 1310
rect 11260 750 11280 1310
rect 11200 730 11280 750
rect 11310 1310 11390 1330
rect 11310 750 11330 1310
rect 11370 750 11390 1310
rect 11310 730 11390 750
rect 11420 1310 11500 1330
rect 11420 750 11440 1310
rect 11480 750 11500 1310
rect 11420 730 11500 750
rect 11530 1310 11610 1330
rect 11530 750 11550 1310
rect 11590 750 11610 1310
rect 11530 730 11610 750
rect 11640 1310 11720 1330
rect 11640 750 11660 1310
rect 11700 750 11720 1310
rect 11640 730 11720 750
rect 11750 1310 11830 1330
rect 11750 750 11770 1310
rect 11810 750 11830 1310
rect 11750 730 11830 750
rect 11860 1310 11940 1330
rect 11860 750 11880 1310
rect 11920 750 11940 1310
rect 11860 730 11940 750
rect 11970 1310 12050 1330
rect 11970 750 11990 1310
rect 12030 750 12050 1310
rect 11970 730 12050 750
rect 12080 1310 12160 1330
rect 12080 750 12100 1310
rect 12140 750 12160 1310
rect 12080 730 12160 750
rect 12190 1310 12270 1330
rect 12190 750 12210 1310
rect 12250 750 12270 1310
rect 12190 730 12270 750
rect 12300 1310 12380 1330
rect 12300 750 12320 1310
rect 12360 750 12380 1310
rect 12300 730 12380 750
rect 12410 1310 12490 1330
rect 12410 750 12430 1310
rect 12470 750 12490 1310
rect 12410 730 12490 750
rect 12520 1310 12600 1330
rect 12520 750 12540 1310
rect 12580 750 12600 1310
rect 12520 730 12600 750
rect 12630 1310 12710 1330
rect 12630 750 12650 1310
rect 12690 750 12710 1310
rect 12630 730 12710 750
rect 12740 1310 12820 1330
rect 12740 750 12760 1310
rect 12800 750 12820 1310
rect 12740 730 12820 750
rect 12850 1310 12930 1330
rect 12850 750 12870 1310
rect 12910 750 12930 1310
rect 12850 730 12930 750
rect 12960 1310 13040 1330
rect 12960 750 12980 1310
rect 13020 750 13040 1310
rect 12960 730 13040 750
rect 13070 1310 13150 1330
rect 13070 750 13090 1310
rect 13130 750 13150 1310
rect 13070 730 13150 750
rect 13180 1310 13250 1330
rect 13180 750 13200 1310
rect 13240 750 13250 1310
rect 13180 730 13250 750
rect 13630 1300 13700 1320
rect 13630 740 13640 1300
rect 13680 740 13700 1300
rect 13630 720 13700 740
rect 13730 1300 13810 1320
rect 13730 740 13750 1300
rect 13790 740 13810 1300
rect 13730 720 13810 740
rect 13840 1300 13920 1320
rect 13840 740 13860 1300
rect 13900 740 13920 1300
rect 13840 720 13920 740
rect 13950 1300 14030 1320
rect 13950 740 13970 1300
rect 14010 740 14030 1300
rect 13950 720 14030 740
rect 14060 1300 14140 1320
rect 14060 740 14080 1300
rect 14120 740 14140 1300
rect 14060 720 14140 740
rect 14170 1300 14250 1320
rect 14170 740 14190 1300
rect 14230 740 14250 1300
rect 14170 720 14250 740
rect 14280 1300 14360 1320
rect 14280 740 14300 1300
rect 14340 740 14360 1300
rect 14280 720 14360 740
rect 14390 1300 14470 1320
rect 14390 740 14410 1300
rect 14450 740 14470 1300
rect 14390 720 14470 740
rect 14500 1300 14580 1320
rect 14500 740 14520 1300
rect 14560 740 14580 1300
rect 14500 720 14580 740
rect 14610 1300 14690 1320
rect 14610 740 14630 1300
rect 14670 740 14690 1300
rect 14610 720 14690 740
rect 14720 1300 14800 1320
rect 14720 740 14740 1300
rect 14780 740 14800 1300
rect 14720 720 14800 740
rect 14830 1300 14910 1320
rect 14830 740 14850 1300
rect 14890 740 14910 1300
rect 14830 720 14910 740
rect 14940 1300 15020 1320
rect 14940 740 14960 1300
rect 15000 740 15020 1300
rect 14940 720 15020 740
rect 15050 1300 15130 1320
rect 15050 740 15070 1300
rect 15110 740 15130 1300
rect 15050 720 15130 740
rect 15160 1300 15240 1320
rect 15160 740 15180 1300
rect 15220 740 15240 1300
rect 15160 720 15240 740
rect 15270 1300 15350 1320
rect 15270 740 15290 1300
rect 15330 740 15350 1300
rect 15270 720 15350 740
rect 15380 1300 15460 1320
rect 15380 740 15400 1300
rect 15440 740 15460 1300
rect 15380 720 15460 740
rect 15490 1300 15570 1320
rect 15490 740 15510 1300
rect 15550 740 15570 1300
rect 15490 720 15570 740
rect 15600 1300 15680 1320
rect 15600 740 15620 1300
rect 15660 740 15680 1300
rect 15600 720 15680 740
rect 15710 1300 15790 1320
rect 15710 740 15730 1300
rect 15770 740 15790 1300
rect 15710 720 15790 740
rect 15820 1300 15900 1320
rect 15820 740 15840 1300
rect 15880 740 15900 1300
rect 15820 720 15900 740
rect 15930 1300 16010 1320
rect 15930 740 15950 1300
rect 15990 740 16010 1300
rect 15930 720 16010 740
rect 16040 1300 16120 1320
rect 16040 740 16060 1300
rect 16100 740 16120 1300
rect 16040 720 16120 740
rect 16150 1300 16230 1320
rect 16150 740 16170 1300
rect 16210 740 16230 1300
rect 16150 720 16230 740
rect 16260 1300 16340 1320
rect 16260 740 16280 1300
rect 16320 740 16340 1300
rect 16260 720 16340 740
rect 16370 1300 16450 1320
rect 16370 740 16390 1300
rect 16430 740 16450 1300
rect 16370 720 16450 740
rect 16480 1300 16560 1320
rect 16480 740 16500 1300
rect 16540 740 16560 1300
rect 16480 720 16560 740
rect 16590 1300 16670 1320
rect 16590 740 16610 1300
rect 16650 740 16670 1300
rect 16590 720 16670 740
rect 16700 1300 16780 1320
rect 16700 740 16720 1300
rect 16760 740 16780 1300
rect 16700 720 16780 740
rect 16810 1300 16890 1320
rect 16810 740 16830 1300
rect 16870 740 16890 1300
rect 16810 720 16890 740
rect 16920 1300 16990 1320
rect 16920 740 16940 1300
rect 16980 740 16990 1300
rect 16920 720 16990 740
<< pdiff >>
rect 23460 43160 23530 43180
rect 21720 42860 21790 42880
rect 21720 42200 21730 42860
rect 21770 42200 21790 42860
rect 21720 42180 21790 42200
rect 21820 42860 21890 42880
rect 21820 42200 21840 42860
rect 21880 42200 21890 42860
rect 21820 42180 21890 42200
rect 21950 42860 22020 42880
rect 21950 42200 21960 42860
rect 22000 42200 22020 42860
rect 21950 42180 22020 42200
rect 22050 42860 22120 42880
rect 22050 42200 22070 42860
rect 22110 42200 22120 42860
rect 22050 42180 22120 42200
rect 22580 42870 22650 42890
rect 22580 42210 22590 42870
rect 22630 42210 22650 42870
rect 22580 42190 22650 42210
rect 22680 42870 22750 42890
rect 22680 42210 22700 42870
rect 22740 42210 22750 42870
rect 22680 42190 22750 42210
rect 22880 42870 22950 42890
rect 22880 42210 22890 42870
rect 22930 42210 22950 42870
rect 22880 42190 22950 42210
rect 22980 42870 23060 42890
rect 22980 42210 23000 42870
rect 23040 42210 23060 42870
rect 22980 42190 23060 42210
rect 23090 42870 23160 42890
rect 23090 42210 23110 42870
rect 23150 42210 23160 42870
rect 23460 42500 23470 43160
rect 23510 42500 23530 43160
rect 23460 42480 23530 42500
rect 23560 43160 23630 43180
rect 23560 42500 23580 43160
rect 23620 42500 23630 43160
rect 23560 42480 23630 42500
rect 23090 42190 23160 42210
rect 2559 41900 2629 41920
rect 2559 41740 2569 41900
rect 2609 41740 2629 41900
rect 2559 41720 2629 41740
rect 2659 41900 2739 41920
rect 2659 41740 2679 41900
rect 2719 41740 2739 41900
rect 2659 41720 2739 41740
rect 2769 41900 2849 41920
rect 2769 41740 2789 41900
rect 2829 41740 2849 41900
rect 2769 41720 2849 41740
rect 2879 41900 2949 41920
rect 2879 41740 2899 41900
rect 2939 41740 2949 41900
rect 2879 41720 2949 41740
rect 3389 41800 3459 41820
rect 2439 41380 2509 41400
rect 2439 41020 2449 41380
rect 2489 41020 2509 41380
rect 2439 41000 2509 41020
rect 2539 41380 2619 41400
rect 2539 41020 2559 41380
rect 2599 41020 2619 41380
rect 2539 41000 2619 41020
rect 2649 41380 2729 41400
rect 2649 41020 2669 41380
rect 2709 41020 2729 41380
rect 2649 41000 2729 41020
rect 2759 41380 2839 41400
rect 2759 41020 2779 41380
rect 2819 41020 2839 41380
rect 2759 41000 2839 41020
rect 2869 41380 2949 41400
rect 2869 41020 2889 41380
rect 2929 41020 2949 41380
rect 2869 41000 2949 41020
rect 2979 41380 3049 41400
rect 2979 41020 2999 41380
rect 3039 41020 3049 41380
rect 3389 41090 3399 41800
rect 3439 41090 3459 41800
rect 3389 41070 3459 41090
rect 3489 41800 3569 41820
rect 3489 41090 3509 41800
rect 3549 41090 3569 41800
rect 3489 41070 3569 41090
rect 3599 41800 3679 41820
rect 3599 41090 3619 41800
rect 3659 41090 3679 41800
rect 3599 41070 3679 41090
rect 3709 41800 3789 41820
rect 3709 41090 3729 41800
rect 3769 41090 3789 41800
rect 3709 41070 3789 41090
rect 3819 41800 3899 41820
rect 3819 41090 3839 41800
rect 3879 41090 3899 41800
rect 3819 41070 3899 41090
rect 3929 41800 4009 41820
rect 3929 41090 3949 41800
rect 3989 41090 4009 41800
rect 3929 41070 4009 41090
rect 4039 41800 4119 41820
rect 4039 41090 4059 41800
rect 4099 41090 4119 41800
rect 4039 41070 4119 41090
rect 4149 41800 4229 41820
rect 4149 41090 4169 41800
rect 4209 41090 4229 41800
rect 4149 41070 4229 41090
rect 4259 41800 4329 41820
rect 5949 41820 6019 41840
rect 4259 41090 4279 41800
rect 4319 41090 4329 41800
rect 4259 41070 4329 41090
rect 4539 41790 4609 41810
rect 4539 41080 4549 41790
rect 4589 41080 4609 41790
rect 2979 41000 3049 41020
rect 4539 41060 4609 41080
rect 4639 41790 4719 41810
rect 4639 41080 4659 41790
rect 4699 41080 4719 41790
rect 4639 41060 4719 41080
rect 4749 41790 4829 41810
rect 4749 41080 4769 41790
rect 4809 41080 4829 41790
rect 4749 41060 4829 41080
rect 4859 41790 4939 41810
rect 4859 41080 4879 41790
rect 4919 41080 4939 41790
rect 4859 41060 4939 41080
rect 4969 41790 5049 41810
rect 4969 41080 4989 41790
rect 5029 41080 5049 41790
rect 4969 41060 5049 41080
rect 5079 41790 5159 41810
rect 5079 41080 5099 41790
rect 5139 41080 5159 41790
rect 5079 41060 5159 41080
rect 5189 41790 5269 41810
rect 5189 41080 5209 41790
rect 5249 41080 5269 41790
rect 5189 41060 5269 41080
rect 5299 41790 5379 41810
rect 5299 41080 5319 41790
rect 5359 41080 5379 41790
rect 5299 41060 5379 41080
rect 5409 41790 5479 41810
rect 5409 41080 5429 41790
rect 5469 41080 5479 41790
rect 5949 41360 5959 41820
rect 5999 41360 6019 41820
rect 5949 41340 6019 41360
rect 6049 41820 6119 41840
rect 6049 41360 6069 41820
rect 6109 41360 6119 41820
rect 6049 41340 6119 41360
rect 6179 41820 6249 41840
rect 6179 41360 6189 41820
rect 6229 41360 6249 41820
rect 6179 41340 6249 41360
rect 6279 41820 6359 41840
rect 6279 41360 6299 41820
rect 6339 41360 6359 41820
rect 6279 41340 6359 41360
rect 6389 41820 6459 41840
rect 6389 41360 6409 41820
rect 6449 41360 6459 41820
rect 6389 41340 6459 41360
rect 6519 41820 6589 41840
rect 6519 41360 6529 41820
rect 6569 41360 6589 41820
rect 6519 41340 6589 41360
rect 6619 41820 6699 41840
rect 6619 41360 6639 41820
rect 6679 41360 6699 41820
rect 6619 41340 6699 41360
rect 6729 41820 6809 41840
rect 6729 41360 6749 41820
rect 6789 41360 6809 41820
rect 6729 41340 6809 41360
rect 6839 41820 6919 41840
rect 6839 41360 6859 41820
rect 6899 41360 6919 41820
rect 6839 41340 6919 41360
rect 6949 41820 7019 41840
rect 6949 41360 6969 41820
rect 7009 41360 7019 41820
rect 6949 41340 7019 41360
rect 7079 41820 7149 41840
rect 7079 41360 7089 41820
rect 7129 41360 7149 41820
rect 7079 41340 7149 41360
rect 7179 41820 7259 41840
rect 7179 41360 7199 41820
rect 7239 41360 7259 41820
rect 7179 41340 7259 41360
rect 7289 41820 7369 41840
rect 7289 41360 7309 41820
rect 7349 41360 7369 41820
rect 7289 41340 7369 41360
rect 7399 41820 7479 41840
rect 7399 41360 7419 41820
rect 7459 41360 7479 41820
rect 7399 41340 7479 41360
rect 7509 41820 7589 41840
rect 7509 41360 7529 41820
rect 7569 41360 7589 41820
rect 7509 41340 7589 41360
rect 7619 41820 7699 41840
rect 7619 41360 7639 41820
rect 7679 41360 7699 41820
rect 7619 41340 7699 41360
rect 7729 41820 7809 41840
rect 7729 41360 7749 41820
rect 7789 41360 7809 41820
rect 7729 41340 7809 41360
rect 7839 41820 7919 41840
rect 7839 41360 7859 41820
rect 7899 41360 7919 41820
rect 7839 41340 7919 41360
rect 7949 41820 8019 41840
rect 7949 41360 7969 41820
rect 8009 41360 8019 41820
rect 7949 41340 8019 41360
rect 8139 41820 8209 41840
rect 8139 41360 8149 41820
rect 8189 41360 8209 41820
rect 8139 41340 8209 41360
rect 8239 41820 8319 41840
rect 8239 41360 8259 41820
rect 8299 41360 8319 41820
rect 8239 41340 8319 41360
rect 8349 41820 8429 41840
rect 8349 41360 8369 41820
rect 8409 41360 8429 41820
rect 8349 41340 8429 41360
rect 8459 41820 8539 41840
rect 8459 41360 8479 41820
rect 8519 41360 8539 41820
rect 8459 41340 8539 41360
rect 8569 41820 8649 41840
rect 8569 41360 8589 41820
rect 8629 41360 8649 41820
rect 8569 41340 8649 41360
rect 8679 41820 8759 41840
rect 8679 41360 8699 41820
rect 8739 41360 8759 41820
rect 8679 41340 8759 41360
rect 8789 41820 8869 41840
rect 8789 41360 8809 41820
rect 8849 41360 8869 41820
rect 8789 41340 8869 41360
rect 8899 41820 8979 41840
rect 8899 41360 8919 41820
rect 8959 41360 8979 41820
rect 8899 41340 8979 41360
rect 9009 41820 9089 41840
rect 9009 41360 9029 41820
rect 9069 41360 9089 41820
rect 9009 41340 9089 41360
rect 9119 41820 9199 41840
rect 9119 41360 9139 41820
rect 9179 41360 9199 41820
rect 9119 41340 9199 41360
rect 9229 41820 9309 41840
rect 9229 41360 9249 41820
rect 9289 41360 9309 41820
rect 9229 41340 9309 41360
rect 9339 41820 9419 41840
rect 9339 41360 9359 41820
rect 9399 41360 9419 41820
rect 9339 41340 9419 41360
rect 9449 41820 9529 41840
rect 9449 41360 9469 41820
rect 9509 41360 9529 41820
rect 9449 41340 9529 41360
rect 9559 41820 9639 41840
rect 9559 41360 9579 41820
rect 9619 41360 9639 41820
rect 9559 41340 9639 41360
rect 9669 41820 9749 41840
rect 9669 41360 9689 41820
rect 9729 41360 9749 41820
rect 9669 41340 9749 41360
rect 9779 41820 9859 41840
rect 9779 41360 9799 41820
rect 9839 41360 9859 41820
rect 9779 41340 9859 41360
rect 9889 41820 9959 41840
rect 9889 41360 9909 41820
rect 9949 41360 9959 41820
rect 9889 41340 9959 41360
rect 5409 41060 5479 41080
rect 3260 40510 3329 40530
rect 3260 39800 3269 40510
rect 3309 39800 3329 40510
rect 3260 39780 3329 39800
rect 3359 40510 3439 40530
rect 3359 39800 3379 40510
rect 3419 39800 3439 40510
rect 3359 39780 3439 39800
rect 3469 40510 3549 40530
rect 3469 39800 3489 40510
rect 3529 39800 3549 40510
rect 3469 39780 3549 39800
rect 3579 40510 3659 40530
rect 3579 39800 3599 40510
rect 3639 39800 3659 40510
rect 3579 39780 3659 39800
rect 3689 40510 3769 40530
rect 3689 39800 3709 40510
rect 3749 39800 3769 40510
rect 3689 39780 3769 39800
rect 3799 40510 3879 40530
rect 3799 39800 3819 40510
rect 3859 39800 3879 40510
rect 3799 39780 3879 39800
rect 3909 40510 3989 40530
rect 3909 39800 3929 40510
rect 3969 39800 3989 40510
rect 3909 39780 3989 39800
rect 4019 40510 4099 40530
rect 4019 39800 4039 40510
rect 4079 39800 4099 40510
rect 4019 39780 4099 39800
rect 4129 40510 4200 40530
rect 4129 39800 4149 40510
rect 4189 39800 4200 40510
rect 4129 39780 4200 39800
rect 4539 40510 4609 40530
rect 4539 39800 4549 40510
rect 4589 39800 4609 40510
rect 4539 39780 4609 39800
rect 4639 40510 4719 40530
rect 4639 39800 4659 40510
rect 4699 39800 4719 40510
rect 4639 39780 4719 39800
rect 4749 40510 4829 40530
rect 4749 39800 4769 40510
rect 4809 39800 4829 40510
rect 4749 39780 4829 39800
rect 4859 40510 4939 40530
rect 4859 39800 4879 40510
rect 4919 39800 4939 40510
rect 4859 39780 4939 39800
rect 4969 40510 5049 40530
rect 4969 39800 4989 40510
rect 5029 39800 5049 40510
rect 4969 39780 5049 39800
rect 5079 40510 5159 40530
rect 5079 39800 5099 40510
rect 5139 39800 5159 40510
rect 5079 39780 5159 39800
rect 5189 40510 5269 40530
rect 5189 39800 5209 40510
rect 5249 39800 5269 40510
rect 5189 39780 5269 39800
rect 5299 40510 5379 40530
rect 5299 39800 5319 40510
rect 5359 39800 5379 40510
rect 5299 39780 5379 39800
rect 5409 40510 5479 40530
rect 5409 39800 5429 40510
rect 5469 39800 5479 40510
rect 6349 40500 6419 40520
rect 6349 40040 6359 40500
rect 6399 40040 6419 40500
rect 6349 40020 6419 40040
rect 6449 40500 6529 40520
rect 6449 40040 6469 40500
rect 6509 40040 6529 40500
rect 6449 40020 6529 40040
rect 6559 40500 6639 40520
rect 6559 40040 6579 40500
rect 6619 40040 6639 40500
rect 6559 40020 6639 40040
rect 6669 40500 6749 40520
rect 6669 40040 6689 40500
rect 6729 40040 6749 40500
rect 6669 40020 6749 40040
rect 6779 40500 6859 40520
rect 6779 40040 6799 40500
rect 6839 40040 6859 40500
rect 6779 40020 6859 40040
rect 6889 40500 6969 40520
rect 6889 40040 6909 40500
rect 6949 40040 6969 40500
rect 6889 40020 6969 40040
rect 6999 40500 7079 40520
rect 6999 40040 7019 40500
rect 7059 40040 7079 40500
rect 6999 40020 7079 40040
rect 7109 40500 7189 40520
rect 7109 40040 7129 40500
rect 7169 40040 7189 40500
rect 7109 40020 7189 40040
rect 7219 40500 7299 40520
rect 7219 40040 7239 40500
rect 7279 40040 7299 40500
rect 7219 40020 7299 40040
rect 7329 40500 7409 40520
rect 7329 40040 7349 40500
rect 7389 40040 7409 40500
rect 7329 40020 7409 40040
rect 7439 40500 7519 40520
rect 7439 40040 7459 40500
rect 7499 40040 7519 40500
rect 7439 40020 7519 40040
rect 7549 40500 7629 40520
rect 7549 40040 7569 40500
rect 7609 40040 7629 40500
rect 7549 40020 7629 40040
rect 7659 40500 7739 40520
rect 7659 40040 7679 40500
rect 7719 40040 7739 40500
rect 7659 40020 7739 40040
rect 7769 40500 7849 40520
rect 7769 40040 7789 40500
rect 7829 40040 7849 40500
rect 7769 40020 7849 40040
rect 7879 40500 7959 40520
rect 7879 40040 7899 40500
rect 7939 40040 7959 40500
rect 7879 40020 7959 40040
rect 7989 40500 8069 40520
rect 7989 40040 8009 40500
rect 8049 40040 8069 40500
rect 7989 40020 8069 40040
rect 8099 40500 8179 40520
rect 8099 40040 8119 40500
rect 8159 40040 8179 40500
rect 8099 40020 8179 40040
rect 8209 40500 8289 40520
rect 8209 40040 8229 40500
rect 8269 40040 8289 40500
rect 8209 40020 8289 40040
rect 8319 40500 8399 40520
rect 8319 40040 8339 40500
rect 8379 40040 8399 40500
rect 8319 40020 8399 40040
rect 8429 40500 8509 40520
rect 8429 40040 8449 40500
rect 8489 40040 8509 40500
rect 8429 40020 8509 40040
rect 8539 40500 8619 40520
rect 8539 40040 8559 40500
rect 8599 40040 8619 40500
rect 8539 40020 8619 40040
rect 8649 40500 8729 40520
rect 8649 40040 8669 40500
rect 8709 40040 8729 40500
rect 8649 40020 8729 40040
rect 8759 40500 8839 40520
rect 8759 40040 8779 40500
rect 8819 40040 8839 40500
rect 8759 40020 8839 40040
rect 8869 40500 8949 40520
rect 8869 40040 8889 40500
rect 8929 40040 8949 40500
rect 8869 40020 8949 40040
rect 8979 40500 9059 40520
rect 8979 40040 8999 40500
rect 9039 40040 9059 40500
rect 8979 40020 9059 40040
rect 9089 40500 9169 40520
rect 9089 40040 9109 40500
rect 9149 40040 9169 40500
rect 9089 40020 9169 40040
rect 9199 40500 9279 40520
rect 9199 40040 9219 40500
rect 9259 40040 9279 40500
rect 9199 40020 9279 40040
rect 9309 40500 9389 40520
rect 9309 40040 9329 40500
rect 9369 40040 9389 40500
rect 9309 40020 9389 40040
rect 9419 40500 9499 40520
rect 9419 40040 9439 40500
rect 9479 40040 9499 40500
rect 9419 40020 9499 40040
rect 9529 40500 9609 40520
rect 9529 40040 9549 40500
rect 9589 40040 9609 40500
rect 9529 40020 9609 40040
rect 9639 40500 9719 40520
rect 9639 40040 9659 40500
rect 9699 40040 9719 40500
rect 9639 40020 9719 40040
rect 9749 40500 9829 40520
rect 9749 40040 9769 40500
rect 9809 40040 9829 40500
rect 9749 40020 9829 40040
rect 9859 40500 9929 40520
rect 9859 40040 9879 40500
rect 9919 40040 9929 40500
rect 9859 40020 9929 40040
rect 5409 39780 5479 39800
rect 5460 34740 5530 34760
rect 3770 34670 3840 34690
rect 3770 33710 3780 34670
rect 3820 33710 3840 34670
rect 3770 33690 3840 33710
rect 3870 34670 3950 34690
rect 3870 33710 3890 34670
rect 3930 33710 3950 34670
rect 3870 33690 3950 33710
rect 3980 34670 4060 34690
rect 3980 33710 4000 34670
rect 4040 33710 4060 34670
rect 3980 33690 4060 33710
rect 4090 34670 4170 34690
rect 4090 33710 4110 34670
rect 4150 33710 4170 34670
rect 4090 33690 4170 33710
rect 4200 34670 4280 34690
rect 4200 33710 4220 34670
rect 4260 33710 4280 34670
rect 4200 33690 4280 33710
rect 4310 34670 4390 34690
rect 4310 33710 4330 34670
rect 4370 33710 4390 34670
rect 4310 33690 4390 33710
rect 4420 34670 4650 34690
rect 4420 33710 4510 34670
rect 4560 33710 4650 34670
rect 4420 33690 4650 33710
rect 4680 34670 4760 34690
rect 4680 33710 4700 34670
rect 4740 33710 4760 34670
rect 4680 33690 4760 33710
rect 4790 34670 4870 34690
rect 4790 33710 4810 34670
rect 4850 33710 4870 34670
rect 4790 33690 4870 33710
rect 4900 34670 4980 34690
rect 4900 33710 4920 34670
rect 4960 33710 4980 34670
rect 4900 33690 4980 33710
rect 5010 34670 5090 34690
rect 5010 33710 5030 34670
rect 5070 33710 5090 34670
rect 5010 33690 5090 33710
rect 5120 34670 5200 34690
rect 5120 33710 5140 34670
rect 5180 33710 5200 34670
rect 5120 33690 5200 33710
rect 5230 34670 5300 34690
rect 5230 33710 5250 34670
rect 5290 33710 5300 34670
rect 5460 33780 5470 34740
rect 5510 33780 5530 34740
rect 5460 33760 5530 33780
rect 5560 34740 5640 34760
rect 5560 33780 5580 34740
rect 5620 33780 5640 34740
rect 5560 33760 5640 33780
rect 5670 34740 5750 34760
rect 5670 33780 5690 34740
rect 5730 33780 5750 34740
rect 5670 33760 5750 33780
rect 5780 34740 5860 34760
rect 5780 33780 5800 34740
rect 5840 33780 5860 34740
rect 5780 33760 5860 33780
rect 5890 34740 5970 34760
rect 5890 33780 5910 34740
rect 5950 33780 5970 34740
rect 5890 33760 5970 33780
rect 6000 34740 6080 34760
rect 6000 33780 6020 34740
rect 6060 33780 6080 34740
rect 6000 33760 6080 33780
rect 6110 34740 6180 34760
rect 6110 33780 6130 34740
rect 6170 33780 6180 34740
rect 6340 34740 6410 34760
rect 6340 34280 6350 34740
rect 6390 34280 6410 34740
rect 6340 34260 6410 34280
rect 6440 34740 6520 34760
rect 6440 34280 6460 34740
rect 6500 34280 6520 34740
rect 6440 34260 6520 34280
rect 6550 34740 6620 34760
rect 19760 36080 19830 36100
rect 17460 36060 17530 36080
rect 15340 35950 15410 35970
rect 15340 35790 15350 35950
rect 15390 35790 15410 35950
rect 15340 35770 15410 35790
rect 15440 35950 15520 35970
rect 15440 35790 15460 35950
rect 15500 35790 15520 35950
rect 15440 35770 15520 35790
rect 15550 35950 15620 35970
rect 15550 35790 15570 35950
rect 15610 35790 15620 35950
rect 15550 35770 15620 35790
rect 17460 35600 17470 36060
rect 17510 35600 17530 36060
rect 17460 35580 17530 35600
rect 17560 36060 17630 36080
rect 17560 35600 17580 36060
rect 17620 35600 17630 36060
rect 17560 35580 17630 35600
rect 17710 36060 17780 36080
rect 17710 35600 17720 36060
rect 17760 35600 17780 36060
rect 17710 35580 17780 35600
rect 17810 36060 17880 36080
rect 17810 35600 17830 36060
rect 17870 35600 17880 36060
rect 17810 35580 17880 35600
rect 18030 36060 18100 36080
rect 18030 35600 18040 36060
rect 18080 35600 18100 36060
rect 18030 35580 18100 35600
rect 18130 36060 18200 36080
rect 18130 35600 18150 36060
rect 18190 35600 18200 36060
rect 18130 35580 18200 35600
rect 18400 36060 18470 36080
rect 18400 35600 18410 36060
rect 18450 35600 18470 36060
rect 18400 35580 18470 35600
rect 18500 36060 18570 36080
rect 18500 35600 18520 36060
rect 18560 35600 18570 36060
rect 18500 35580 18570 35600
rect 18650 36060 18720 36080
rect 18650 35600 18660 36060
rect 18700 35600 18720 36060
rect 18650 35580 18720 35600
rect 18750 36060 18820 36080
rect 18750 35600 18770 36060
rect 18810 35600 18820 36060
rect 18750 35580 18820 35600
rect 18970 36060 19040 36080
rect 18970 35600 18980 36060
rect 19020 35600 19040 36060
rect 18970 35580 19040 35600
rect 19070 36060 19140 36080
rect 19070 35600 19090 36060
rect 19130 35600 19140 36060
rect 19070 35580 19140 35600
rect 19300 35990 19370 36010
rect 6550 34280 6570 34740
rect 6610 34280 6620 34740
rect 6550 34260 6620 34280
rect 6700 34250 6770 34750
rect 6800 34730 6880 34750
rect 6800 34270 6820 34730
rect 6860 34270 6880 34730
rect 6800 34250 6880 34270
rect 6910 34730 7030 34750
rect 6910 34270 6950 34730
rect 6990 34270 7030 34730
rect 6910 34250 7030 34270
rect 7060 34730 7140 34750
rect 7060 34270 7080 34730
rect 7120 34270 7140 34730
rect 7060 34250 7140 34270
rect 7170 34250 7240 34750
rect 7300 34730 7370 34750
rect 7300 34270 7310 34730
rect 7350 34270 7370 34730
rect 7300 34250 7370 34270
rect 7400 34730 7480 34750
rect 7400 34270 7420 34730
rect 7460 34270 7480 34730
rect 7400 34250 7480 34270
rect 7510 34730 7580 34750
rect 7510 34270 7530 34730
rect 7570 34270 7580 34730
rect 7510 34250 7580 34270
rect 7680 34730 7750 34750
rect 7680 34270 7690 34730
rect 7730 34270 7750 34730
rect 7680 34250 7750 34270
rect 7780 34730 7860 34750
rect 7780 34270 7800 34730
rect 7840 34270 7860 34730
rect 7780 34250 7860 34270
rect 7890 34730 7960 34750
rect 7890 34270 7910 34730
rect 7950 34270 7960 34730
rect 7890 34250 7960 34270
rect 8060 34730 8130 34750
rect 8060 34270 8070 34730
rect 8110 34270 8130 34730
rect 8060 34250 8130 34270
rect 8160 34730 8240 34750
rect 8160 34270 8180 34730
rect 8220 34270 8240 34730
rect 8160 34250 8240 34270
rect 8270 34730 8340 34750
rect 8270 34270 8290 34730
rect 8330 34270 8340 34730
rect 8270 34250 8340 34270
rect 8440 34730 8510 34750
rect 8440 34270 8450 34730
rect 8490 34270 8510 34730
rect 8440 34250 8510 34270
rect 8540 34730 8620 34750
rect 8540 34270 8560 34730
rect 8600 34270 8620 34730
rect 8540 34250 8620 34270
rect 8650 34730 8720 34750
rect 8650 34270 8670 34730
rect 8710 34270 8720 34730
rect 8650 34250 8720 34270
rect 8780 34250 8850 34750
rect 8880 34730 8960 34750
rect 8880 34270 8900 34730
rect 8940 34270 8960 34730
rect 8880 34250 8960 34270
rect 8990 34730 9110 34750
rect 8990 34270 9030 34730
rect 9070 34270 9110 34730
rect 8990 34250 9110 34270
rect 9140 34730 9220 34750
rect 9140 34270 9160 34730
rect 9200 34270 9220 34730
rect 9140 34250 9220 34270
rect 9250 34250 9320 34750
rect 9380 34730 9450 34750
rect 9380 34270 9390 34730
rect 9430 34270 9450 34730
rect 9380 34250 9450 34270
rect 9480 34730 9560 34750
rect 9480 34270 9500 34730
rect 9540 34270 9560 34730
rect 9480 34250 9560 34270
rect 9590 34730 9660 34750
rect 9590 34270 9610 34730
rect 9650 34270 9660 34730
rect 9590 34250 9660 34270
rect 9760 34730 9830 34750
rect 9760 34270 9770 34730
rect 9810 34270 9830 34730
rect 9760 34250 9830 34270
rect 9860 34730 9940 34750
rect 9860 34270 9880 34730
rect 9920 34270 9940 34730
rect 9860 34250 9940 34270
rect 9970 34730 10040 34750
rect 9970 34270 9990 34730
rect 10030 34270 10040 34730
rect 9970 34250 10040 34270
rect 10140 34730 10210 34750
rect 10140 34270 10150 34730
rect 10190 34270 10210 34730
rect 10140 34250 10210 34270
rect 10240 34730 10320 34750
rect 10240 34270 10260 34730
rect 10300 34270 10320 34730
rect 10240 34250 10320 34270
rect 10350 34730 10420 34750
rect 10350 34270 10370 34730
rect 10410 34270 10420 34730
rect 10350 34250 10420 34270
rect 10520 34730 10590 34750
rect 10520 34270 10530 34730
rect 10570 34270 10590 34730
rect 10520 34250 10590 34270
rect 10620 34730 10700 34750
rect 10620 34270 10640 34730
rect 10680 34270 10700 34730
rect 10620 34250 10700 34270
rect 10730 34730 10800 34750
rect 10730 34270 10750 34730
rect 10790 34270 10800 34730
rect 19300 35030 19310 35990
rect 19350 35030 19370 35990
rect 19300 35010 19370 35030
rect 19400 35990 19470 36010
rect 19400 35030 19420 35990
rect 19460 35030 19470 35990
rect 19760 35620 19770 36080
rect 19810 35620 19830 36080
rect 19760 35600 19830 35620
rect 19860 36080 19930 36100
rect 19860 35620 19880 36080
rect 19920 35620 19930 36080
rect 19860 35600 19930 35620
rect 20010 36080 20080 36100
rect 20010 35620 20020 36080
rect 20060 35620 20080 36080
rect 20010 35600 20080 35620
rect 20110 36080 20180 36100
rect 24720 36080 24790 36100
rect 20110 35620 20130 36080
rect 20170 35620 20180 36080
rect 22420 36060 22490 36080
rect 20110 35600 20180 35620
rect 21030 35990 21100 36010
rect 19400 35010 19470 35030
rect 21030 35030 21040 35990
rect 21080 35030 21100 35990
rect 21030 35010 21100 35030
rect 21130 35990 21200 36010
rect 21130 35030 21150 35990
rect 21190 35030 21200 35990
rect 22420 35600 22430 36060
rect 22470 35600 22490 36060
rect 22420 35580 22490 35600
rect 22520 36060 22590 36080
rect 22520 35600 22540 36060
rect 22580 35600 22590 36060
rect 22520 35580 22590 35600
rect 22670 36060 22740 36080
rect 22670 35600 22680 36060
rect 22720 35600 22740 36060
rect 22670 35580 22740 35600
rect 22770 36060 22840 36080
rect 22770 35600 22790 36060
rect 22830 35600 22840 36060
rect 22770 35580 22840 35600
rect 22990 36060 23060 36080
rect 22990 35600 23000 36060
rect 23040 35600 23060 36060
rect 22990 35580 23060 35600
rect 23090 36060 23160 36080
rect 23090 35600 23110 36060
rect 23150 35600 23160 36060
rect 23090 35580 23160 35600
rect 23360 36060 23430 36080
rect 23360 35600 23370 36060
rect 23410 35600 23430 36060
rect 23360 35580 23430 35600
rect 23460 36060 23530 36080
rect 23460 35600 23480 36060
rect 23520 35600 23530 36060
rect 23460 35580 23530 35600
rect 23610 36060 23680 36080
rect 23610 35600 23620 36060
rect 23660 35600 23680 36060
rect 23610 35580 23680 35600
rect 23710 36060 23780 36080
rect 23710 35600 23730 36060
rect 23770 35600 23780 36060
rect 23710 35580 23780 35600
rect 23930 36060 24000 36080
rect 23930 35600 23940 36060
rect 23980 35600 24000 36060
rect 23930 35580 24000 35600
rect 24030 36060 24100 36080
rect 24030 35600 24050 36060
rect 24090 35600 24100 36060
rect 24030 35580 24100 35600
rect 24260 35990 24330 36010
rect 21130 35010 21200 35030
rect 24260 35030 24270 35990
rect 24310 35030 24330 35990
rect 24260 35010 24330 35030
rect 24360 35990 24430 36010
rect 24360 35030 24380 35990
rect 24420 35030 24430 35990
rect 24720 35620 24730 36080
rect 24770 35620 24790 36080
rect 24720 35600 24790 35620
rect 24820 36080 24890 36100
rect 24820 35620 24840 36080
rect 24880 35620 24890 36080
rect 24820 35600 24890 35620
rect 24970 36080 25040 36100
rect 24970 35620 24980 36080
rect 25020 35620 25040 36080
rect 24970 35600 25040 35620
rect 25070 36080 25140 36100
rect 25070 35620 25090 36080
rect 25130 35620 25140 36080
rect 25070 35600 25140 35620
rect 24360 35010 24430 35030
rect 10730 34250 10800 34270
rect 6110 33760 6180 33780
rect 5230 33690 5300 33710
rect 13888 32220 13958 32240
rect 13888 32060 13898 32220
rect 13938 32060 13958 32220
rect 13888 32040 13958 32060
rect 13988 32220 14068 32240
rect 13988 32060 14008 32220
rect 14048 32060 14068 32220
rect 13988 32040 14068 32060
rect 14098 32220 14178 32240
rect 14098 32060 14118 32220
rect 14158 32060 14178 32220
rect 14098 32040 14178 32060
rect 14208 32220 14278 32240
rect 14208 32060 14228 32220
rect 14268 32060 14278 32220
rect 14208 32040 14278 32060
rect 17460 32000 17530 32020
rect 17460 31540 17470 32000
rect 17510 31540 17530 32000
rect 17460 31520 17530 31540
rect 17560 32000 17630 32020
rect 17560 31540 17580 32000
rect 17620 31540 17630 32000
rect 17560 31520 17630 31540
rect 17710 32000 17780 32020
rect 17710 31540 17720 32000
rect 17760 31540 17780 32000
rect 17710 31520 17780 31540
rect 17810 32000 17880 32020
rect 17810 31540 17830 32000
rect 17870 31540 17880 32000
rect 17810 31520 17880 31540
rect 18030 32000 18100 32020
rect 18030 31540 18040 32000
rect 18080 31540 18100 32000
rect 18030 31520 18100 31540
rect 18130 32000 18200 32020
rect 18130 31540 18150 32000
rect 18190 31540 18200 32000
rect 18130 31520 18200 31540
rect 18400 32000 18470 32020
rect 18400 31540 18410 32000
rect 18450 31540 18470 32000
rect 18400 31520 18470 31540
rect 18500 32000 18570 32020
rect 18500 31540 18520 32000
rect 18560 31540 18570 32000
rect 18500 31520 18570 31540
rect 18650 32000 18720 32020
rect 18650 31540 18660 32000
rect 18700 31540 18720 32000
rect 18650 31520 18720 31540
rect 18750 32000 18820 32020
rect 18750 31540 18770 32000
rect 18810 31540 18820 32000
rect 18750 31520 18820 31540
rect 18970 32000 19040 32020
rect 18970 31540 18980 32000
rect 19020 31540 19040 32000
rect 18970 31520 19040 31540
rect 19070 32000 19140 32020
rect 19070 31540 19090 32000
rect 19130 31540 19140 32000
rect 20020 32000 20090 32020
rect 19070 31520 19140 31540
rect 19300 31930 19370 31950
rect 6400 30590 6470 30610
rect 3860 30490 3930 30510
rect 2170 30420 2240 30440
rect 2170 29460 2180 30420
rect 2220 29460 2240 30420
rect 2170 29440 2240 29460
rect 2270 30420 2350 30440
rect 2270 29460 2290 30420
rect 2330 29460 2350 30420
rect 2270 29440 2350 29460
rect 2380 30420 2460 30440
rect 2380 29460 2400 30420
rect 2440 29460 2460 30420
rect 2380 29440 2460 29460
rect 2490 30420 2570 30440
rect 2490 29460 2510 30420
rect 2550 29460 2570 30420
rect 2490 29440 2570 29460
rect 2600 30420 2680 30440
rect 2600 29460 2620 30420
rect 2660 29460 2680 30420
rect 2600 29440 2680 29460
rect 2710 30420 2790 30440
rect 2710 29460 2730 30420
rect 2770 29460 2790 30420
rect 2710 29440 2790 29460
rect 2820 30420 3050 30440
rect 2820 29460 2910 30420
rect 2960 29460 3050 30420
rect 2820 29440 3050 29460
rect 3080 30420 3160 30440
rect 3080 29460 3100 30420
rect 3140 29460 3160 30420
rect 3080 29440 3160 29460
rect 3190 30420 3270 30440
rect 3190 29460 3210 30420
rect 3250 29460 3270 30420
rect 3190 29440 3270 29460
rect 3300 30420 3380 30440
rect 3300 29460 3320 30420
rect 3360 29460 3380 30420
rect 3300 29440 3380 29460
rect 3410 30420 3490 30440
rect 3410 29460 3430 30420
rect 3470 29460 3490 30420
rect 3410 29440 3490 29460
rect 3520 30420 3600 30440
rect 3520 29460 3540 30420
rect 3580 29460 3600 30420
rect 3520 29440 3600 29460
rect 3630 30420 3700 30440
rect 3630 29460 3650 30420
rect 3690 29460 3700 30420
rect 3860 29530 3870 30490
rect 3910 29530 3930 30490
rect 3860 29510 3930 29530
rect 3960 30490 4040 30510
rect 3960 29530 3980 30490
rect 4020 29530 4040 30490
rect 3960 29510 4040 29530
rect 4070 30490 4150 30510
rect 4070 29530 4090 30490
rect 4130 29530 4150 30490
rect 4070 29510 4150 29530
rect 4180 30490 4260 30510
rect 4180 29530 4200 30490
rect 4240 29530 4260 30490
rect 4180 29510 4260 29530
rect 4290 30490 4370 30510
rect 4290 29530 4310 30490
rect 4350 29530 4370 30490
rect 4290 29510 4370 29530
rect 4400 30490 4480 30510
rect 4400 29530 4420 30490
rect 4460 29530 4480 30490
rect 4400 29510 4480 29530
rect 4510 30490 4580 30510
rect 4510 29530 4530 30490
rect 4570 29530 4580 30490
rect 4510 29510 4580 29530
rect 4720 30490 4790 30510
rect 4720 29530 4730 30490
rect 4770 29530 4790 30490
rect 4720 29510 4790 29530
rect 4820 30490 4900 30510
rect 4820 29530 4840 30490
rect 4880 29530 4900 30490
rect 4820 29510 4900 29530
rect 4930 30490 5010 30510
rect 4930 29530 4950 30490
rect 4990 29530 5010 30490
rect 4930 29510 5010 29530
rect 5040 30490 5120 30510
rect 5040 29530 5060 30490
rect 5100 29530 5120 30490
rect 5040 29510 5120 29530
rect 5150 30490 5230 30510
rect 5150 29530 5170 30490
rect 5210 29530 5230 30490
rect 5150 29510 5230 29530
rect 5260 30490 5340 30510
rect 5260 29530 5280 30490
rect 5320 29530 5340 30490
rect 5260 29510 5340 29530
rect 5370 30490 5440 30510
rect 5370 29530 5390 30490
rect 5430 29530 5440 30490
rect 5370 29510 5440 29530
rect 5580 30490 5650 30510
rect 5580 29530 5590 30490
rect 5630 29530 5650 30490
rect 5580 29510 5650 29530
rect 5680 30490 5760 30510
rect 5680 29530 5700 30490
rect 5740 29530 5760 30490
rect 5680 29510 5760 29530
rect 5790 30490 5870 30510
rect 5790 29530 5810 30490
rect 5850 29530 5870 30490
rect 5790 29510 5870 29530
rect 5900 30490 5980 30510
rect 5900 29530 5920 30490
rect 5960 29530 5980 30490
rect 5900 29510 5980 29530
rect 6010 30490 6090 30510
rect 6010 29530 6030 30490
rect 6070 29530 6090 30490
rect 6010 29510 6090 29530
rect 6120 30490 6200 30510
rect 6120 29530 6140 30490
rect 6180 29530 6200 30490
rect 6120 29510 6200 29530
rect 6230 30490 6300 30510
rect 6230 29530 6250 30490
rect 6290 29530 6300 30490
rect 6400 30130 6410 30590
rect 6450 30130 6470 30590
rect 6400 30110 6470 30130
rect 6500 30590 6580 30610
rect 6500 30130 6520 30590
rect 6560 30130 6580 30590
rect 6500 30110 6580 30130
rect 6610 30590 6680 30610
rect 6610 30130 6630 30590
rect 6670 30130 6680 30590
rect 6610 30110 6680 30130
rect 6760 30100 6830 30600
rect 6860 30580 6940 30600
rect 6860 30120 6880 30580
rect 6920 30120 6940 30580
rect 6860 30100 6940 30120
rect 6970 30580 7090 30600
rect 6970 30120 7010 30580
rect 7050 30120 7090 30580
rect 6970 30100 7090 30120
rect 7120 30580 7200 30600
rect 7120 30120 7140 30580
rect 7180 30120 7200 30580
rect 7120 30100 7200 30120
rect 7230 30100 7300 30600
rect 7360 30580 7430 30600
rect 7360 30120 7370 30580
rect 7410 30120 7430 30580
rect 7360 30100 7430 30120
rect 7460 30580 7540 30600
rect 7460 30120 7480 30580
rect 7520 30120 7540 30580
rect 7460 30100 7540 30120
rect 7570 30580 7640 30600
rect 7570 30120 7590 30580
rect 7630 30120 7640 30580
rect 7570 30100 7640 30120
rect 7740 30580 7810 30600
rect 7740 30120 7750 30580
rect 7790 30120 7810 30580
rect 7740 30100 7810 30120
rect 7840 30580 7920 30600
rect 7840 30120 7860 30580
rect 7900 30120 7920 30580
rect 7840 30100 7920 30120
rect 7950 30580 8020 30600
rect 7950 30120 7970 30580
rect 8010 30120 8020 30580
rect 7950 30100 8020 30120
rect 8120 30580 8190 30600
rect 8120 30120 8130 30580
rect 8170 30120 8190 30580
rect 8120 30100 8190 30120
rect 8220 30580 8300 30600
rect 8220 30120 8240 30580
rect 8280 30120 8300 30580
rect 8220 30100 8300 30120
rect 8330 30580 8400 30600
rect 8330 30120 8350 30580
rect 8390 30120 8400 30580
rect 8330 30100 8400 30120
rect 8500 30580 8570 30600
rect 8500 30120 8510 30580
rect 8550 30120 8570 30580
rect 8500 30100 8570 30120
rect 8600 30580 8680 30600
rect 8600 30120 8620 30580
rect 8660 30120 8680 30580
rect 8600 30100 8680 30120
rect 8710 30580 8780 30600
rect 8710 30120 8730 30580
rect 8770 30120 8780 30580
rect 8710 30100 8780 30120
rect 8840 30100 8910 30600
rect 8940 30580 9020 30600
rect 8940 30120 8960 30580
rect 9000 30120 9020 30580
rect 8940 30100 9020 30120
rect 9050 30580 9170 30600
rect 9050 30120 9090 30580
rect 9130 30120 9170 30580
rect 9050 30100 9170 30120
rect 9200 30580 9280 30600
rect 9200 30120 9220 30580
rect 9260 30120 9280 30580
rect 9200 30100 9280 30120
rect 9310 30100 9380 30600
rect 9440 30580 9510 30600
rect 9440 30120 9450 30580
rect 9490 30120 9510 30580
rect 9440 30100 9510 30120
rect 9540 30580 9620 30600
rect 9540 30120 9560 30580
rect 9600 30120 9620 30580
rect 9540 30100 9620 30120
rect 9650 30580 9720 30600
rect 9650 30120 9670 30580
rect 9710 30120 9720 30580
rect 9650 30100 9720 30120
rect 9820 30580 9890 30600
rect 9820 30120 9830 30580
rect 9870 30120 9890 30580
rect 9820 30100 9890 30120
rect 9920 30580 10000 30600
rect 9920 30120 9940 30580
rect 9980 30120 10000 30580
rect 9920 30100 10000 30120
rect 10030 30580 10100 30600
rect 10030 30120 10050 30580
rect 10090 30120 10100 30580
rect 10030 30100 10100 30120
rect 10200 30580 10270 30600
rect 10200 30120 10210 30580
rect 10250 30120 10270 30580
rect 10200 30100 10270 30120
rect 10300 30580 10380 30600
rect 10300 30120 10320 30580
rect 10360 30120 10380 30580
rect 10300 30100 10380 30120
rect 10410 30580 10480 30600
rect 10410 30120 10430 30580
rect 10470 30120 10480 30580
rect 10410 30100 10480 30120
rect 10580 30580 10650 30600
rect 10580 30120 10590 30580
rect 10630 30120 10650 30580
rect 10580 30100 10650 30120
rect 10680 30580 10760 30600
rect 10680 30120 10700 30580
rect 10740 30120 10760 30580
rect 10680 30100 10760 30120
rect 10790 30580 10860 30600
rect 10790 30120 10810 30580
rect 10850 30120 10860 30580
rect 10790 30100 10860 30120
rect 10960 30580 11030 30600
rect 10960 30120 10970 30580
rect 11010 30120 11030 30580
rect 10960 30100 11030 30120
rect 11060 30580 11140 30600
rect 11060 30120 11080 30580
rect 11120 30120 11140 30580
rect 11060 30100 11140 30120
rect 11170 30580 11240 30600
rect 11170 30120 11190 30580
rect 11230 30120 11240 30580
rect 19300 30970 19310 31930
rect 19350 30970 19370 31930
rect 19300 30950 19370 30970
rect 19400 31930 19470 31950
rect 19400 30970 19420 31930
rect 19460 30970 19470 31930
rect 19400 30950 19470 30970
rect 19560 31930 19630 31950
rect 19560 30970 19570 31930
rect 19610 30970 19630 31930
rect 19560 30950 19630 30970
rect 19660 31930 19730 31950
rect 19660 30970 19680 31930
rect 19720 30970 19730 31930
rect 20020 31540 20030 32000
rect 20070 31540 20090 32000
rect 20020 31520 20090 31540
rect 20120 32000 20190 32020
rect 20120 31540 20140 32000
rect 20180 31540 20190 32000
rect 20120 31520 20190 31540
rect 20270 32000 20340 32020
rect 20270 31540 20280 32000
rect 20320 31540 20340 32000
rect 20270 31520 20340 31540
rect 20370 32000 20440 32020
rect 24980 32010 25050 32030
rect 20370 31540 20390 32000
rect 20430 31540 20440 32000
rect 22480 31990 22550 32010
rect 20370 31520 20440 31540
rect 21090 31930 21160 31950
rect 19660 30950 19730 30970
rect 21090 30970 21100 31930
rect 21140 30970 21160 31930
rect 21090 30950 21160 30970
rect 21190 31930 21260 31950
rect 21190 30970 21210 31930
rect 21250 30970 21260 31930
rect 22480 31530 22490 31990
rect 22530 31530 22550 31990
rect 22480 31510 22550 31530
rect 22580 31990 22650 32010
rect 22580 31530 22600 31990
rect 22640 31530 22650 31990
rect 22580 31510 22650 31530
rect 22730 31990 22800 32010
rect 22730 31530 22740 31990
rect 22780 31530 22800 31990
rect 22730 31510 22800 31530
rect 22830 31990 22900 32010
rect 22830 31530 22850 31990
rect 22890 31530 22900 31990
rect 22830 31510 22900 31530
rect 23050 31990 23120 32010
rect 23050 31530 23060 31990
rect 23100 31530 23120 31990
rect 23050 31510 23120 31530
rect 23150 31990 23220 32010
rect 23150 31530 23170 31990
rect 23210 31530 23220 31990
rect 23150 31510 23220 31530
rect 23420 31990 23490 32010
rect 23420 31530 23430 31990
rect 23470 31530 23490 31990
rect 23420 31510 23490 31530
rect 23520 31990 23590 32010
rect 23520 31530 23540 31990
rect 23580 31530 23590 31990
rect 23520 31510 23590 31530
rect 23670 31990 23740 32010
rect 23670 31530 23680 31990
rect 23720 31530 23740 31990
rect 23670 31510 23740 31530
rect 23770 31990 23840 32010
rect 23770 31530 23790 31990
rect 23830 31530 23840 31990
rect 23770 31510 23840 31530
rect 23990 31990 24060 32010
rect 23990 31530 24000 31990
rect 24040 31530 24060 31990
rect 23990 31510 24060 31530
rect 24090 31990 24160 32010
rect 24090 31530 24110 31990
rect 24150 31530 24160 31990
rect 24090 31510 24160 31530
rect 24320 31920 24390 31940
rect 21190 30950 21260 30970
rect 24320 30960 24330 31920
rect 24370 30960 24390 31920
rect 24320 30940 24390 30960
rect 24420 31920 24490 31940
rect 24420 30960 24440 31920
rect 24480 30960 24490 31920
rect 24420 30940 24490 30960
rect 24580 31920 24650 31940
rect 24580 30960 24590 31920
rect 24630 30960 24650 31920
rect 24580 30940 24650 30960
rect 24680 31920 24750 31940
rect 24680 30960 24700 31920
rect 24740 30960 24750 31920
rect 24980 31550 24990 32010
rect 25030 31550 25050 32010
rect 24980 31530 25050 31550
rect 25080 32010 25150 32030
rect 25080 31550 25100 32010
rect 25140 31550 25150 32010
rect 25080 31530 25150 31550
rect 25230 32010 25300 32030
rect 25230 31550 25240 32010
rect 25280 31550 25300 32010
rect 25230 31530 25300 31550
rect 25330 32010 25400 32030
rect 25330 31550 25350 32010
rect 25390 31550 25400 32010
rect 25330 31530 25400 31550
rect 24680 30940 24750 30960
rect 11170 30100 11240 30120
rect 6230 29510 6300 29530
rect 3630 29440 3700 29460
rect 7320 26470 7390 26490
rect 7320 26010 7330 26470
rect 7370 26010 7390 26470
rect 7320 25990 7390 26010
rect 7420 26470 7500 26490
rect 7420 26010 7440 26470
rect 7480 26010 7500 26470
rect 7420 25990 7500 26010
rect 7530 26470 7600 26490
rect 7530 26010 7550 26470
rect 7590 26010 7600 26470
rect 7530 25990 7600 26010
rect 7850 26470 7920 26490
rect 7850 26010 7860 26470
rect 7900 26010 7920 26470
rect 7850 25990 7920 26010
rect 7950 26470 8030 26490
rect 7950 26010 7970 26470
rect 8010 26010 8030 26470
rect 7950 25990 8030 26010
rect 8060 26470 8130 26490
rect 8060 26010 8080 26470
rect 8120 26010 8130 26470
rect 8060 25990 8130 26010
rect 8480 26480 8550 26500
rect 8480 26020 8490 26480
rect 8530 26020 8550 26480
rect 8480 26000 8550 26020
rect 8580 26480 8700 26500
rect 8580 26020 8620 26480
rect 8660 26020 8700 26480
rect 8580 26000 8700 26020
rect 8730 26480 8800 26500
rect 8730 26020 8750 26480
rect 8790 26020 8800 26480
rect 8730 26000 8800 26020
rect 8860 26480 8930 26500
rect 8860 26020 8870 26480
rect 8910 26020 8930 26480
rect 8860 26000 8930 26020
rect 8960 26480 9030 26500
rect 8960 26020 8980 26480
rect 9020 26020 9030 26480
rect 8960 26000 9030 26020
rect 9220 26480 9290 26500
rect 9220 26020 9230 26480
rect 9270 26020 9290 26480
rect 9220 26000 9290 26020
rect 9320 26480 9400 26500
rect 9320 26020 9340 26480
rect 9380 26020 9400 26480
rect 9320 26000 9400 26020
rect 9430 26480 9500 26500
rect 9430 26020 9450 26480
rect 9490 26020 9500 26480
rect 9430 26000 9500 26020
rect 9560 26000 9630 26500
rect 9660 26480 9740 26500
rect 9660 26020 9680 26480
rect 9720 26020 9740 26480
rect 9660 26000 9740 26020
rect 9770 26480 9890 26500
rect 9770 26020 9810 26480
rect 9850 26020 9890 26480
rect 9770 26000 9890 26020
rect 9920 26480 10000 26500
rect 9920 26020 9940 26480
rect 9980 26020 10000 26480
rect 9920 26000 10000 26020
rect 10030 26000 10100 26500
rect 10160 26480 10230 26500
rect 10160 26020 10170 26480
rect 10210 26020 10230 26480
rect 10160 26000 10230 26020
rect 10260 26480 10340 26500
rect 10260 26020 10280 26480
rect 10320 26020 10340 26480
rect 10260 26000 10340 26020
rect 10370 26480 10440 26500
rect 10370 26020 10390 26480
rect 10430 26020 10440 26480
rect 10370 26000 10440 26020
rect 10550 26000 10620 26500
rect 10650 26480 10730 26500
rect 10650 26020 10670 26480
rect 10710 26020 10730 26480
rect 10650 26000 10730 26020
rect 10760 26480 10880 26500
rect 10760 26020 10800 26480
rect 10840 26020 10880 26480
rect 10760 26000 10880 26020
rect 10910 26480 10990 26500
rect 10910 26020 10930 26480
rect 10970 26020 10990 26480
rect 10910 26000 10990 26020
rect 11020 26000 11090 26500
rect 11150 26480 11220 26500
rect 11150 26020 11160 26480
rect 11200 26020 11220 26480
rect 11150 26000 11220 26020
rect 11250 26480 11330 26500
rect 11250 26020 11270 26480
rect 11310 26020 11330 26480
rect 11250 26000 11330 26020
rect 11360 26480 11430 26500
rect 11360 26020 11380 26480
rect 11420 26020 11430 26480
rect 11360 26000 11430 26020
rect 11550 26000 11620 26500
rect 11650 26480 11730 26500
rect 11650 26020 11670 26480
rect 11710 26020 11730 26480
rect 11650 26000 11730 26020
rect 11760 26480 11880 26500
rect 11760 26020 11800 26480
rect 11840 26020 11880 26480
rect 11760 26000 11880 26020
rect 11910 26480 11990 26500
rect 11910 26020 11930 26480
rect 11970 26020 11990 26480
rect 11910 26000 11990 26020
rect 12020 26000 12090 26500
rect 12150 26480 12220 26500
rect 12150 26020 12160 26480
rect 12200 26020 12220 26480
rect 12150 26000 12220 26020
rect 12250 26480 12330 26500
rect 12250 26020 12270 26480
rect 12310 26020 12330 26480
rect 12250 26000 12330 26020
rect 12360 26480 12430 26500
rect 12360 26020 12380 26480
rect 12420 26020 12430 26480
rect 12360 26000 12430 26020
rect 12530 26480 12600 26500
rect 12530 26020 12540 26480
rect 12580 26020 12600 26480
rect 12530 26000 12600 26020
rect 12630 26480 12710 26500
rect 12630 26020 12650 26480
rect 12690 26020 12710 26480
rect 12630 26000 12710 26020
rect 12740 26480 12810 26500
rect 12740 26020 12760 26480
rect 12800 26020 12810 26480
rect 12740 26000 12810 26020
rect 12880 26480 12950 26500
rect 12880 26020 12890 26480
rect 12930 26020 12950 26480
rect 12880 26000 12950 26020
rect 12980 26480 13050 26500
rect 12980 26020 13000 26480
rect 13040 26020 13050 26480
rect 12980 26000 13050 26020
rect 13110 26480 13180 26500
rect 13110 26020 13120 26480
rect 13160 26020 13180 26480
rect 13110 26000 13180 26020
rect 13210 26480 13290 26500
rect 13210 26020 13230 26480
rect 13270 26020 13290 26480
rect 13210 26000 13290 26020
rect 13320 26480 13390 26500
rect 13320 26020 13340 26480
rect 13380 26020 13390 26480
rect 13320 26000 13390 26020
rect 13450 26480 13520 26500
rect 13450 26020 13460 26480
rect 13500 26020 13520 26480
rect 13450 26000 13520 26020
rect 13550 26480 13630 26500
rect 13550 26020 13570 26480
rect 13610 26020 13630 26480
rect 13550 26000 13630 26020
rect 13660 26480 13740 26500
rect 13660 26020 13680 26480
rect 13720 26020 13740 26480
rect 13660 26000 13740 26020
rect 13770 26480 13850 26500
rect 13770 26020 13790 26480
rect 13830 26020 13850 26480
rect 13770 26000 13850 26020
rect 13880 26480 13950 26500
rect 13880 26020 13900 26480
rect 13940 26020 13950 26480
rect 13880 26000 13950 26020
rect 14010 26480 14080 26500
rect 14010 26020 14020 26480
rect 14060 26020 14080 26480
rect 14010 26000 14080 26020
rect 14110 26480 14190 26500
rect 14110 26020 14130 26480
rect 14170 26020 14190 26480
rect 14110 26000 14190 26020
rect 14220 26480 14300 26500
rect 14220 26020 14240 26480
rect 14280 26020 14300 26480
rect 14220 26000 14300 26020
rect 14330 26480 14410 26500
rect 14330 26020 14350 26480
rect 14390 26020 14410 26480
rect 14330 26000 14410 26020
rect 14440 26480 14520 26500
rect 14440 26020 14460 26480
rect 14500 26020 14520 26480
rect 14440 26000 14520 26020
rect 14550 26480 14630 26500
rect 14550 26020 14570 26480
rect 14610 26020 14630 26480
rect 14550 26000 14630 26020
rect 14660 26480 14740 26500
rect 14660 26020 14680 26480
rect 14720 26020 14740 26480
rect 14660 26000 14740 26020
rect 14770 26480 14850 26500
rect 14770 26020 14790 26480
rect 14830 26020 14850 26480
rect 14770 26000 14850 26020
rect 14880 26480 14950 26500
rect 14880 26020 14900 26480
rect 14940 26020 14950 26480
rect 14880 26000 14950 26020
rect 15070 26480 15140 26500
rect 15070 26020 15080 26480
rect 15120 26020 15140 26480
rect 15070 26000 15140 26020
rect 15170 26480 15250 26500
rect 15170 26020 15190 26480
rect 15230 26020 15250 26480
rect 15170 26000 15250 26020
rect 15280 26480 15360 26500
rect 15280 26020 15300 26480
rect 15340 26020 15360 26480
rect 15280 26000 15360 26020
rect 15390 26480 15470 26500
rect 15390 26020 15410 26480
rect 15450 26020 15470 26480
rect 15390 26000 15470 26020
rect 15500 26480 15580 26500
rect 15500 26020 15520 26480
rect 15560 26020 15580 26480
rect 15500 26000 15580 26020
rect 15610 26480 15690 26500
rect 15610 26020 15630 26480
rect 15670 26020 15690 26480
rect 15610 26000 15690 26020
rect 15720 26480 15800 26500
rect 15720 26020 15740 26480
rect 15780 26020 15800 26480
rect 15720 26000 15800 26020
rect 15830 26480 15910 26500
rect 15830 26020 15850 26480
rect 15890 26020 15910 26480
rect 15830 26000 15910 26020
rect 15940 26480 16020 26500
rect 15940 26020 15960 26480
rect 16000 26020 16020 26480
rect 15940 26000 16020 26020
rect 16050 26480 16130 26500
rect 16050 26020 16070 26480
rect 16110 26020 16130 26480
rect 16050 26000 16130 26020
rect 16160 26480 16240 26500
rect 16160 26020 16180 26480
rect 16220 26020 16240 26480
rect 16160 26000 16240 26020
rect 16270 26480 16350 26500
rect 16270 26020 16290 26480
rect 16330 26020 16350 26480
rect 16270 26000 16350 26020
rect 16380 26480 16460 26500
rect 16380 26020 16400 26480
rect 16440 26020 16460 26480
rect 16380 26000 16460 26020
rect 16490 26480 16570 26500
rect 16490 26020 16510 26480
rect 16550 26020 16570 26480
rect 16490 26000 16570 26020
rect 16600 26480 16680 26500
rect 16600 26020 16620 26480
rect 16660 26020 16680 26480
rect 16600 26000 16680 26020
rect 16710 26480 16790 26500
rect 16710 26020 16730 26480
rect 16770 26020 16790 26480
rect 16710 26000 16790 26020
rect 16820 26480 16890 26500
rect 16820 26020 16840 26480
rect 16880 26020 16890 26480
rect 16820 26000 16890 26020
rect 17020 26480 17090 26500
rect 17020 26020 17030 26480
rect 17070 26020 17090 26480
rect 17020 26000 17090 26020
rect 17120 26480 17200 26500
rect 17120 26020 17140 26480
rect 17180 26020 17200 26480
rect 17120 26000 17200 26020
rect 17230 26480 17310 26500
rect 17230 26020 17250 26480
rect 17290 26020 17310 26480
rect 17230 26000 17310 26020
rect 17340 26480 17420 26500
rect 17340 26020 17360 26480
rect 17400 26020 17420 26480
rect 17340 26000 17420 26020
rect 17450 26480 17530 26500
rect 17450 26020 17470 26480
rect 17510 26020 17530 26480
rect 17450 26000 17530 26020
rect 17560 26480 17640 26500
rect 17560 26020 17580 26480
rect 17620 26020 17640 26480
rect 17560 26000 17640 26020
rect 17670 26480 17750 26500
rect 17670 26020 17690 26480
rect 17730 26020 17750 26480
rect 17670 26000 17750 26020
rect 17780 26480 17860 26500
rect 17780 26020 17800 26480
rect 17840 26020 17860 26480
rect 17780 26000 17860 26020
rect 17890 26480 17970 26500
rect 17890 26020 17910 26480
rect 17950 26020 17970 26480
rect 17890 26000 17970 26020
rect 18000 26480 18080 26500
rect 18000 26020 18020 26480
rect 18060 26020 18080 26480
rect 18000 26000 18080 26020
rect 18110 26480 18190 26500
rect 18110 26020 18130 26480
rect 18170 26020 18190 26480
rect 18110 26000 18190 26020
rect 18220 26480 18300 26500
rect 18220 26020 18240 26480
rect 18280 26020 18300 26480
rect 18220 26000 18300 26020
rect 18330 26480 18410 26500
rect 18330 26020 18350 26480
rect 18390 26020 18410 26480
rect 18330 26000 18410 26020
rect 18440 26480 18520 26500
rect 18440 26020 18460 26480
rect 18500 26020 18520 26480
rect 18440 26000 18520 26020
rect 18550 26480 18630 26500
rect 18550 26020 18570 26480
rect 18610 26020 18630 26480
rect 18550 26000 18630 26020
rect 18660 26480 18740 26500
rect 18660 26020 18680 26480
rect 18720 26020 18740 26480
rect 18660 26000 18740 26020
rect 18770 26480 18850 26500
rect 18770 26020 18790 26480
rect 18830 26020 18850 26480
rect 18770 26000 18850 26020
rect 18880 26480 18960 26500
rect 18880 26020 18900 26480
rect 18940 26020 18960 26480
rect 18880 26000 18960 26020
rect 18990 26480 19070 26500
rect 18990 26020 19010 26480
rect 19050 26020 19070 26480
rect 18990 26000 19070 26020
rect 19100 26480 19180 26500
rect 19100 26020 19120 26480
rect 19160 26020 19180 26480
rect 19100 26000 19180 26020
rect 19210 26480 19290 26500
rect 19210 26020 19230 26480
rect 19270 26020 19290 26480
rect 19210 26000 19290 26020
rect 19320 26480 19400 26500
rect 19320 26020 19340 26480
rect 19380 26020 19400 26480
rect 19320 26000 19400 26020
rect 19430 26480 19510 26500
rect 19430 26020 19450 26480
rect 19490 26020 19510 26480
rect 19430 26000 19510 26020
rect 19540 26480 19620 26500
rect 19540 26020 19560 26480
rect 19600 26020 19620 26480
rect 19540 26000 19620 26020
rect 19650 26480 19730 26500
rect 19650 26020 19670 26480
rect 19710 26020 19730 26480
rect 19650 26000 19730 26020
rect 19760 26480 19840 26500
rect 19760 26020 19780 26480
rect 19820 26020 19840 26480
rect 19760 26000 19840 26020
rect 19870 26480 19950 26500
rect 19870 26020 19890 26480
rect 19930 26020 19950 26480
rect 19870 26000 19950 26020
rect 19980 26480 20060 26500
rect 19980 26020 20000 26480
rect 20040 26020 20060 26480
rect 19980 26000 20060 26020
rect 20090 26480 20170 26500
rect 20090 26020 20110 26480
rect 20150 26020 20170 26480
rect 20090 26000 20170 26020
rect 20200 26480 20280 26500
rect 20200 26020 20220 26480
rect 20260 26020 20280 26480
rect 20200 26000 20280 26020
rect 20310 26480 20390 26500
rect 20310 26020 20330 26480
rect 20370 26020 20390 26480
rect 20310 26000 20390 26020
rect 20420 26480 20500 26500
rect 20420 26020 20440 26480
rect 20480 26020 20500 26480
rect 20420 26000 20500 26020
rect 20530 26480 20600 26500
rect 20530 26020 20550 26480
rect 20590 26020 20600 26480
rect 20530 26000 20600 26020
rect 7360 21080 7430 21580
rect 7460 21560 7540 21580
rect 7460 21100 7480 21560
rect 7520 21100 7540 21560
rect 7460 21080 7540 21100
rect 7570 21560 7690 21580
rect 7570 21100 7610 21560
rect 7650 21100 7690 21560
rect 7570 21080 7690 21100
rect 7720 21560 7800 21580
rect 7720 21100 7740 21560
rect 7780 21100 7800 21560
rect 7720 21080 7800 21100
rect 7830 21080 7900 21580
rect 7960 21560 8030 21580
rect 7960 21100 7970 21560
rect 8010 21100 8030 21560
rect 7960 21080 8030 21100
rect 8060 21560 8140 21580
rect 8060 21100 8080 21560
rect 8120 21100 8140 21560
rect 8060 21080 8140 21100
rect 8170 21560 8240 21580
rect 8170 21100 8190 21560
rect 8230 21100 8240 21560
rect 8170 21080 8240 21100
rect 8480 21550 8550 21570
rect 8480 21090 8490 21550
rect 8530 21090 8550 21550
rect 8480 21070 8550 21090
rect 8580 21550 8700 21570
rect 8580 21090 8620 21550
rect 8660 21090 8700 21550
rect 8580 21070 8700 21090
rect 8730 21550 8800 21570
rect 8730 21090 8750 21550
rect 8790 21090 8800 21550
rect 8730 21070 8800 21090
rect 8860 21550 8930 21570
rect 8860 21090 8870 21550
rect 8910 21090 8930 21550
rect 8860 21070 8930 21090
rect 8960 21550 9030 21570
rect 8960 21090 8980 21550
rect 9020 21090 9030 21550
rect 8960 21070 9030 21090
rect 9220 21550 9290 21570
rect 9220 21090 9230 21550
rect 9270 21090 9290 21550
rect 9220 21070 9290 21090
rect 9320 21550 9400 21570
rect 9320 21090 9340 21550
rect 9380 21090 9400 21550
rect 9320 21070 9400 21090
rect 9430 21550 9500 21570
rect 9430 21090 9450 21550
rect 9490 21090 9500 21550
rect 9430 21070 9500 21090
rect 9560 21070 9630 21570
rect 9660 21550 9740 21570
rect 9660 21090 9680 21550
rect 9720 21090 9740 21550
rect 9660 21070 9740 21090
rect 9770 21550 9890 21570
rect 9770 21090 9810 21550
rect 9850 21090 9890 21550
rect 9770 21070 9890 21090
rect 9920 21550 10000 21570
rect 9920 21090 9940 21550
rect 9980 21090 10000 21550
rect 9920 21070 10000 21090
rect 10030 21070 10100 21570
rect 10160 21550 10230 21570
rect 10160 21090 10170 21550
rect 10210 21090 10230 21550
rect 10160 21070 10230 21090
rect 10260 21550 10340 21570
rect 10260 21090 10280 21550
rect 10320 21090 10340 21550
rect 10260 21070 10340 21090
rect 10370 21550 10440 21570
rect 10370 21090 10390 21550
rect 10430 21090 10440 21550
rect 10370 21070 10440 21090
rect 10550 21070 10620 21570
rect 10650 21550 10730 21570
rect 10650 21090 10670 21550
rect 10710 21090 10730 21550
rect 10650 21070 10730 21090
rect 10760 21550 10880 21570
rect 10760 21090 10800 21550
rect 10840 21090 10880 21550
rect 10760 21070 10880 21090
rect 10910 21550 10990 21570
rect 10910 21090 10930 21550
rect 10970 21090 10990 21550
rect 10910 21070 10990 21090
rect 11020 21070 11090 21570
rect 11150 21550 11220 21570
rect 11150 21090 11160 21550
rect 11200 21090 11220 21550
rect 11150 21070 11220 21090
rect 11250 21550 11330 21570
rect 11250 21090 11270 21550
rect 11310 21090 11330 21550
rect 11250 21070 11330 21090
rect 11360 21550 11430 21570
rect 11360 21090 11380 21550
rect 11420 21090 11430 21550
rect 11360 21070 11430 21090
rect 11550 21070 11620 21570
rect 11650 21550 11730 21570
rect 11650 21090 11670 21550
rect 11710 21090 11730 21550
rect 11650 21070 11730 21090
rect 11760 21550 11880 21570
rect 11760 21090 11800 21550
rect 11840 21090 11880 21550
rect 11760 21070 11880 21090
rect 11910 21550 11990 21570
rect 11910 21090 11930 21550
rect 11970 21090 11990 21550
rect 11910 21070 11990 21090
rect 12020 21070 12090 21570
rect 12150 21550 12220 21570
rect 12150 21090 12160 21550
rect 12200 21090 12220 21550
rect 12150 21070 12220 21090
rect 12250 21550 12330 21570
rect 12250 21090 12270 21550
rect 12310 21090 12330 21550
rect 12250 21070 12330 21090
rect 12360 21550 12430 21570
rect 12360 21090 12380 21550
rect 12420 21090 12430 21550
rect 12360 21070 12430 21090
rect 12530 21550 12600 21570
rect 12530 21090 12540 21550
rect 12580 21090 12600 21550
rect 12530 21070 12600 21090
rect 12630 21550 12710 21570
rect 12630 21090 12650 21550
rect 12690 21090 12710 21550
rect 12630 21070 12710 21090
rect 12740 21550 12810 21570
rect 12740 21090 12760 21550
rect 12800 21090 12810 21550
rect 12740 21070 12810 21090
rect 12880 21550 12950 21570
rect 12880 21090 12890 21550
rect 12930 21090 12950 21550
rect 12880 21070 12950 21090
rect 12980 21550 13050 21570
rect 12980 21090 13000 21550
rect 13040 21090 13050 21550
rect 12980 21070 13050 21090
rect 13110 21550 13180 21570
rect 13110 21090 13120 21550
rect 13160 21090 13180 21550
rect 13110 21070 13180 21090
rect 13210 21550 13290 21570
rect 13210 21090 13230 21550
rect 13270 21090 13290 21550
rect 13210 21070 13290 21090
rect 13320 21550 13390 21570
rect 13320 21090 13340 21550
rect 13380 21090 13390 21550
rect 13320 21070 13390 21090
rect 13450 21550 13520 21570
rect 13450 21090 13460 21550
rect 13500 21090 13520 21550
rect 13450 21070 13520 21090
rect 13550 21550 13630 21570
rect 13550 21090 13570 21550
rect 13610 21090 13630 21550
rect 13550 21070 13630 21090
rect 13660 21550 13740 21570
rect 13660 21090 13680 21550
rect 13720 21090 13740 21550
rect 13660 21070 13740 21090
rect 13770 21550 13850 21570
rect 13770 21090 13790 21550
rect 13830 21090 13850 21550
rect 13770 21070 13850 21090
rect 13880 21550 13950 21570
rect 13880 21090 13900 21550
rect 13940 21090 13950 21550
rect 13880 21070 13950 21090
rect 14010 21550 14080 21570
rect 14010 21090 14020 21550
rect 14060 21090 14080 21550
rect 14010 21070 14080 21090
rect 14110 21550 14190 21570
rect 14110 21090 14130 21550
rect 14170 21090 14190 21550
rect 14110 21070 14190 21090
rect 14220 21550 14300 21570
rect 14220 21090 14240 21550
rect 14280 21090 14300 21550
rect 14220 21070 14300 21090
rect 14330 21550 14410 21570
rect 14330 21090 14350 21550
rect 14390 21090 14410 21550
rect 14330 21070 14410 21090
rect 14440 21550 14520 21570
rect 14440 21090 14460 21550
rect 14500 21090 14520 21550
rect 14440 21070 14520 21090
rect 14550 21550 14630 21570
rect 14550 21090 14570 21550
rect 14610 21090 14630 21550
rect 14550 21070 14630 21090
rect 14660 21550 14740 21570
rect 14660 21090 14680 21550
rect 14720 21090 14740 21550
rect 14660 21070 14740 21090
rect 14770 21550 14850 21570
rect 14770 21090 14790 21550
rect 14830 21090 14850 21550
rect 14770 21070 14850 21090
rect 14880 21550 14950 21570
rect 14880 21090 14900 21550
rect 14940 21090 14950 21550
rect 14880 21070 14950 21090
rect 15070 21550 15140 21570
rect 15070 21090 15080 21550
rect 15120 21090 15140 21550
rect 15070 21070 15140 21090
rect 15170 21550 15250 21570
rect 15170 21090 15190 21550
rect 15230 21090 15250 21550
rect 15170 21070 15250 21090
rect 15280 21550 15360 21570
rect 15280 21090 15300 21550
rect 15340 21090 15360 21550
rect 15280 21070 15360 21090
rect 15390 21550 15470 21570
rect 15390 21090 15410 21550
rect 15450 21090 15470 21550
rect 15390 21070 15470 21090
rect 15500 21550 15580 21570
rect 15500 21090 15520 21550
rect 15560 21090 15580 21550
rect 15500 21070 15580 21090
rect 15610 21550 15690 21570
rect 15610 21090 15630 21550
rect 15670 21090 15690 21550
rect 15610 21070 15690 21090
rect 15720 21550 15800 21570
rect 15720 21090 15740 21550
rect 15780 21090 15800 21550
rect 15720 21070 15800 21090
rect 15830 21550 15910 21570
rect 15830 21090 15850 21550
rect 15890 21090 15910 21550
rect 15830 21070 15910 21090
rect 15940 21550 16020 21570
rect 15940 21090 15960 21550
rect 16000 21090 16020 21550
rect 15940 21070 16020 21090
rect 16050 21550 16130 21570
rect 16050 21090 16070 21550
rect 16110 21090 16130 21550
rect 16050 21070 16130 21090
rect 16160 21550 16240 21570
rect 16160 21090 16180 21550
rect 16220 21090 16240 21550
rect 16160 21070 16240 21090
rect 16270 21550 16350 21570
rect 16270 21090 16290 21550
rect 16330 21090 16350 21550
rect 16270 21070 16350 21090
rect 16380 21550 16460 21570
rect 16380 21090 16400 21550
rect 16440 21090 16460 21550
rect 16380 21070 16460 21090
rect 16490 21550 16570 21570
rect 16490 21090 16510 21550
rect 16550 21090 16570 21550
rect 16490 21070 16570 21090
rect 16600 21550 16680 21570
rect 16600 21090 16620 21550
rect 16660 21090 16680 21550
rect 16600 21070 16680 21090
rect 16710 21550 16790 21570
rect 16710 21090 16730 21550
rect 16770 21090 16790 21550
rect 16710 21070 16790 21090
rect 16820 21550 16890 21570
rect 16820 21090 16840 21550
rect 16880 21090 16890 21550
rect 16820 21070 16890 21090
rect 17020 21550 17090 21570
rect 17020 21090 17030 21550
rect 17070 21090 17090 21550
rect 17020 21070 17090 21090
rect 17120 21550 17200 21570
rect 17120 21090 17140 21550
rect 17180 21090 17200 21550
rect 17120 21070 17200 21090
rect 17230 21550 17310 21570
rect 17230 21090 17250 21550
rect 17290 21090 17310 21550
rect 17230 21070 17310 21090
rect 17340 21550 17420 21570
rect 17340 21090 17360 21550
rect 17400 21090 17420 21550
rect 17340 21070 17420 21090
rect 17450 21550 17530 21570
rect 17450 21090 17470 21550
rect 17510 21090 17530 21550
rect 17450 21070 17530 21090
rect 17560 21550 17640 21570
rect 17560 21090 17580 21550
rect 17620 21090 17640 21550
rect 17560 21070 17640 21090
rect 17670 21550 17750 21570
rect 17670 21090 17690 21550
rect 17730 21090 17750 21550
rect 17670 21070 17750 21090
rect 17780 21550 17860 21570
rect 17780 21090 17800 21550
rect 17840 21090 17860 21550
rect 17780 21070 17860 21090
rect 17890 21550 17970 21570
rect 17890 21090 17910 21550
rect 17950 21090 17970 21550
rect 17890 21070 17970 21090
rect 18000 21550 18080 21570
rect 18000 21090 18020 21550
rect 18060 21090 18080 21550
rect 18000 21070 18080 21090
rect 18110 21550 18190 21570
rect 18110 21090 18130 21550
rect 18170 21090 18190 21550
rect 18110 21070 18190 21090
rect 18220 21550 18300 21570
rect 18220 21090 18240 21550
rect 18280 21090 18300 21550
rect 18220 21070 18300 21090
rect 18330 21550 18410 21570
rect 18330 21090 18350 21550
rect 18390 21090 18410 21550
rect 18330 21070 18410 21090
rect 18440 21550 18520 21570
rect 18440 21090 18460 21550
rect 18500 21090 18520 21550
rect 18440 21070 18520 21090
rect 18550 21550 18630 21570
rect 18550 21090 18570 21550
rect 18610 21090 18630 21550
rect 18550 21070 18630 21090
rect 18660 21550 18740 21570
rect 18660 21090 18680 21550
rect 18720 21090 18740 21550
rect 18660 21070 18740 21090
rect 18770 21550 18850 21570
rect 18770 21090 18790 21550
rect 18830 21090 18850 21550
rect 18770 21070 18850 21090
rect 18880 21550 18960 21570
rect 18880 21090 18900 21550
rect 18940 21090 18960 21550
rect 18880 21070 18960 21090
rect 18990 21550 19070 21570
rect 18990 21090 19010 21550
rect 19050 21090 19070 21550
rect 18990 21070 19070 21090
rect 19100 21550 19180 21570
rect 19100 21090 19120 21550
rect 19160 21090 19180 21550
rect 19100 21070 19180 21090
rect 19210 21550 19290 21570
rect 19210 21090 19230 21550
rect 19270 21090 19290 21550
rect 19210 21070 19290 21090
rect 19320 21550 19400 21570
rect 19320 21090 19340 21550
rect 19380 21090 19400 21550
rect 19320 21070 19400 21090
rect 19430 21550 19510 21570
rect 19430 21090 19450 21550
rect 19490 21090 19510 21550
rect 19430 21070 19510 21090
rect 19540 21550 19620 21570
rect 19540 21090 19560 21550
rect 19600 21090 19620 21550
rect 19540 21070 19620 21090
rect 19650 21550 19730 21570
rect 19650 21090 19670 21550
rect 19710 21090 19730 21550
rect 19650 21070 19730 21090
rect 19760 21550 19840 21570
rect 19760 21090 19780 21550
rect 19820 21090 19840 21550
rect 19760 21070 19840 21090
rect 19870 21550 19950 21570
rect 19870 21090 19890 21550
rect 19930 21090 19950 21550
rect 19870 21070 19950 21090
rect 19980 21550 20060 21570
rect 19980 21090 20000 21550
rect 20040 21090 20060 21550
rect 19980 21070 20060 21090
rect 20090 21550 20170 21570
rect 20090 21090 20110 21550
rect 20150 21090 20170 21550
rect 20090 21070 20170 21090
rect 20200 21550 20280 21570
rect 20200 21090 20220 21550
rect 20260 21090 20280 21550
rect 20200 21070 20280 21090
rect 20310 21550 20390 21570
rect 20310 21090 20330 21550
rect 20370 21090 20390 21550
rect 20310 21070 20390 21090
rect 20420 21550 20500 21570
rect 20420 21090 20440 21550
rect 20480 21090 20500 21550
rect 20420 21070 20500 21090
rect 20530 21550 20600 21570
rect 20530 21090 20550 21550
rect 20590 21090 20600 21550
rect 20530 21070 20600 21090
rect 7280 19360 7350 20360
rect 7380 20340 7460 20360
rect 7380 19380 7400 20340
rect 7440 19380 7460 20340
rect 7380 19360 7460 19380
rect 7490 19360 7610 20360
rect 7640 20340 7720 20360
rect 7640 19380 7660 20340
rect 7700 19380 7720 20340
rect 7640 19360 7720 19380
rect 7750 19360 7820 20360
rect 7950 20340 8020 20360
rect 7950 19880 7960 20340
rect 8000 19880 8020 20340
rect 7950 19860 8020 19880
rect 8050 20340 8130 20360
rect 8050 19880 8070 20340
rect 8110 19880 8130 20340
rect 8050 19860 8130 19880
rect 8160 20340 8230 20360
rect 8160 19880 8180 20340
rect 8220 19880 8230 20340
rect 8160 19860 8230 19880
rect 8480 19890 8550 19910
rect 8480 19430 8490 19890
rect 8530 19430 8550 19890
rect 8480 19410 8550 19430
rect 8580 19890 8700 19910
rect 8580 19430 8620 19890
rect 8660 19430 8700 19890
rect 8580 19410 8700 19430
rect 8730 19890 8800 19910
rect 8730 19430 8750 19890
rect 8790 19430 8800 19890
rect 8730 19410 8800 19430
rect 8860 19890 8930 19910
rect 8860 19430 8870 19890
rect 8910 19430 8930 19890
rect 8860 19410 8930 19430
rect 8960 19890 9030 19910
rect 8960 19430 8980 19890
rect 9020 19430 9030 19890
rect 8960 19410 9030 19430
rect 9220 19890 9290 19910
rect 9220 19430 9230 19890
rect 9270 19430 9290 19890
rect 9220 19410 9290 19430
rect 9320 19890 9400 19910
rect 9320 19430 9340 19890
rect 9380 19430 9400 19890
rect 9320 19410 9400 19430
rect 9430 19890 9500 19910
rect 9430 19430 9450 19890
rect 9490 19430 9500 19890
rect 9430 19410 9500 19430
rect 9560 19410 9630 19910
rect 9660 19890 9740 19910
rect 9660 19430 9680 19890
rect 9720 19430 9740 19890
rect 9660 19410 9740 19430
rect 9770 19890 9890 19910
rect 9770 19430 9810 19890
rect 9850 19430 9890 19890
rect 9770 19410 9890 19430
rect 9920 19890 10000 19910
rect 9920 19430 9940 19890
rect 9980 19430 10000 19890
rect 9920 19410 10000 19430
rect 10030 19410 10100 19910
rect 10160 19890 10230 19910
rect 10160 19430 10170 19890
rect 10210 19430 10230 19890
rect 10160 19410 10230 19430
rect 10260 19890 10340 19910
rect 10260 19430 10280 19890
rect 10320 19430 10340 19890
rect 10260 19410 10340 19430
rect 10370 19890 10440 19910
rect 10370 19430 10390 19890
rect 10430 19430 10440 19890
rect 10370 19410 10440 19430
rect 10550 19410 10620 19910
rect 10650 19890 10730 19910
rect 10650 19430 10670 19890
rect 10710 19430 10730 19890
rect 10650 19410 10730 19430
rect 10760 19890 10880 19910
rect 10760 19430 10800 19890
rect 10840 19430 10880 19890
rect 10760 19410 10880 19430
rect 10910 19890 10990 19910
rect 10910 19430 10930 19890
rect 10970 19430 10990 19890
rect 10910 19410 10990 19430
rect 11020 19410 11090 19910
rect 11150 19890 11220 19910
rect 11150 19430 11160 19890
rect 11200 19430 11220 19890
rect 11150 19410 11220 19430
rect 11250 19890 11330 19910
rect 11250 19430 11270 19890
rect 11310 19430 11330 19890
rect 11250 19410 11330 19430
rect 11360 19890 11430 19910
rect 11360 19430 11380 19890
rect 11420 19430 11430 19890
rect 11360 19410 11430 19430
rect 11550 19410 11620 19910
rect 11650 19890 11730 19910
rect 11650 19430 11670 19890
rect 11710 19430 11730 19890
rect 11650 19410 11730 19430
rect 11760 19890 11880 19910
rect 11760 19430 11800 19890
rect 11840 19430 11880 19890
rect 11760 19410 11880 19430
rect 11910 19890 11990 19910
rect 11910 19430 11930 19890
rect 11970 19430 11990 19890
rect 11910 19410 11990 19430
rect 12020 19410 12090 19910
rect 12150 19890 12220 19910
rect 12150 19430 12160 19890
rect 12200 19430 12220 19890
rect 12150 19410 12220 19430
rect 12250 19890 12330 19910
rect 12250 19430 12270 19890
rect 12310 19430 12330 19890
rect 12250 19410 12330 19430
rect 12360 19890 12430 19910
rect 12360 19430 12380 19890
rect 12420 19430 12430 19890
rect 12360 19410 12430 19430
rect 12530 19890 12600 19910
rect 12530 19430 12540 19890
rect 12580 19430 12600 19890
rect 12530 19410 12600 19430
rect 12630 19890 12710 19910
rect 12630 19430 12650 19890
rect 12690 19430 12710 19890
rect 12630 19410 12710 19430
rect 12740 19890 12810 19910
rect 12740 19430 12760 19890
rect 12800 19430 12810 19890
rect 12740 19410 12810 19430
rect 12880 19890 12950 19910
rect 12880 19430 12890 19890
rect 12930 19430 12950 19890
rect 12880 19410 12950 19430
rect 12980 19890 13050 19910
rect 12980 19430 13000 19890
rect 13040 19430 13050 19890
rect 12980 19410 13050 19430
rect 13110 19890 13180 19910
rect 13110 19430 13120 19890
rect 13160 19430 13180 19890
rect 13110 19410 13180 19430
rect 13210 19890 13290 19910
rect 13210 19430 13230 19890
rect 13270 19430 13290 19890
rect 13210 19410 13290 19430
rect 13320 19890 13390 19910
rect 13320 19430 13340 19890
rect 13380 19430 13390 19890
rect 13320 19410 13390 19430
rect 13450 19890 13520 19910
rect 13450 19430 13460 19890
rect 13500 19430 13520 19890
rect 13450 19410 13520 19430
rect 13550 19890 13630 19910
rect 13550 19430 13570 19890
rect 13610 19430 13630 19890
rect 13550 19410 13630 19430
rect 13660 19890 13740 19910
rect 13660 19430 13680 19890
rect 13720 19430 13740 19890
rect 13660 19410 13740 19430
rect 13770 19890 13850 19910
rect 13770 19430 13790 19890
rect 13830 19430 13850 19890
rect 13770 19410 13850 19430
rect 13880 19890 13950 19910
rect 13880 19430 13900 19890
rect 13940 19430 13950 19890
rect 13880 19410 13950 19430
rect 14010 19890 14080 19910
rect 14010 19430 14020 19890
rect 14060 19430 14080 19890
rect 14010 19410 14080 19430
rect 14110 19890 14190 19910
rect 14110 19430 14130 19890
rect 14170 19430 14190 19890
rect 14110 19410 14190 19430
rect 14220 19890 14300 19910
rect 14220 19430 14240 19890
rect 14280 19430 14300 19890
rect 14220 19410 14300 19430
rect 14330 19890 14410 19910
rect 14330 19430 14350 19890
rect 14390 19430 14410 19890
rect 14330 19410 14410 19430
rect 14440 19890 14520 19910
rect 14440 19430 14460 19890
rect 14500 19430 14520 19890
rect 14440 19410 14520 19430
rect 14550 19890 14630 19910
rect 14550 19430 14570 19890
rect 14610 19430 14630 19890
rect 14550 19410 14630 19430
rect 14660 19890 14740 19910
rect 14660 19430 14680 19890
rect 14720 19430 14740 19890
rect 14660 19410 14740 19430
rect 14770 19890 14850 19910
rect 14770 19430 14790 19890
rect 14830 19430 14850 19890
rect 14770 19410 14850 19430
rect 14880 19890 14950 19910
rect 14880 19430 14900 19890
rect 14940 19430 14950 19890
rect 14880 19410 14950 19430
rect 15070 19890 15140 19910
rect 15070 19430 15080 19890
rect 15120 19430 15140 19890
rect 15070 19410 15140 19430
rect 15170 19890 15250 19910
rect 15170 19430 15190 19890
rect 15230 19430 15250 19890
rect 15170 19410 15250 19430
rect 15280 19890 15360 19910
rect 15280 19430 15300 19890
rect 15340 19430 15360 19890
rect 15280 19410 15360 19430
rect 15390 19890 15470 19910
rect 15390 19430 15410 19890
rect 15450 19430 15470 19890
rect 15390 19410 15470 19430
rect 15500 19890 15580 19910
rect 15500 19430 15520 19890
rect 15560 19430 15580 19890
rect 15500 19410 15580 19430
rect 15610 19890 15690 19910
rect 15610 19430 15630 19890
rect 15670 19430 15690 19890
rect 15610 19410 15690 19430
rect 15720 19890 15800 19910
rect 15720 19430 15740 19890
rect 15780 19430 15800 19890
rect 15720 19410 15800 19430
rect 15830 19890 15910 19910
rect 15830 19430 15850 19890
rect 15890 19430 15910 19890
rect 15830 19410 15910 19430
rect 15940 19890 16020 19910
rect 15940 19430 15960 19890
rect 16000 19430 16020 19890
rect 15940 19410 16020 19430
rect 16050 19890 16130 19910
rect 16050 19430 16070 19890
rect 16110 19430 16130 19890
rect 16050 19410 16130 19430
rect 16160 19890 16240 19910
rect 16160 19430 16180 19890
rect 16220 19430 16240 19890
rect 16160 19410 16240 19430
rect 16270 19890 16350 19910
rect 16270 19430 16290 19890
rect 16330 19430 16350 19890
rect 16270 19410 16350 19430
rect 16380 19890 16460 19910
rect 16380 19430 16400 19890
rect 16440 19430 16460 19890
rect 16380 19410 16460 19430
rect 16490 19890 16570 19910
rect 16490 19430 16510 19890
rect 16550 19430 16570 19890
rect 16490 19410 16570 19430
rect 16600 19890 16680 19910
rect 16600 19430 16620 19890
rect 16660 19430 16680 19890
rect 16600 19410 16680 19430
rect 16710 19890 16790 19910
rect 16710 19430 16730 19890
rect 16770 19430 16790 19890
rect 16710 19410 16790 19430
rect 16820 19890 16890 19910
rect 16820 19430 16840 19890
rect 16880 19430 16890 19890
rect 16820 19410 16890 19430
rect 17020 19890 17090 19910
rect 17020 19430 17030 19890
rect 17070 19430 17090 19890
rect 17020 19410 17090 19430
rect 17120 19890 17200 19910
rect 17120 19430 17140 19890
rect 17180 19430 17200 19890
rect 17120 19410 17200 19430
rect 17230 19890 17310 19910
rect 17230 19430 17250 19890
rect 17290 19430 17310 19890
rect 17230 19410 17310 19430
rect 17340 19890 17420 19910
rect 17340 19430 17360 19890
rect 17400 19430 17420 19890
rect 17340 19410 17420 19430
rect 17450 19890 17530 19910
rect 17450 19430 17470 19890
rect 17510 19430 17530 19890
rect 17450 19410 17530 19430
rect 17560 19890 17640 19910
rect 17560 19430 17580 19890
rect 17620 19430 17640 19890
rect 17560 19410 17640 19430
rect 17670 19890 17750 19910
rect 17670 19430 17690 19890
rect 17730 19430 17750 19890
rect 17670 19410 17750 19430
rect 17780 19890 17860 19910
rect 17780 19430 17800 19890
rect 17840 19430 17860 19890
rect 17780 19410 17860 19430
rect 17890 19890 17970 19910
rect 17890 19430 17910 19890
rect 17950 19430 17970 19890
rect 17890 19410 17970 19430
rect 18000 19890 18080 19910
rect 18000 19430 18020 19890
rect 18060 19430 18080 19890
rect 18000 19410 18080 19430
rect 18110 19890 18190 19910
rect 18110 19430 18130 19890
rect 18170 19430 18190 19890
rect 18110 19410 18190 19430
rect 18220 19890 18300 19910
rect 18220 19430 18240 19890
rect 18280 19430 18300 19890
rect 18220 19410 18300 19430
rect 18330 19890 18410 19910
rect 18330 19430 18350 19890
rect 18390 19430 18410 19890
rect 18330 19410 18410 19430
rect 18440 19890 18520 19910
rect 18440 19430 18460 19890
rect 18500 19430 18520 19890
rect 18440 19410 18520 19430
rect 18550 19890 18630 19910
rect 18550 19430 18570 19890
rect 18610 19430 18630 19890
rect 18550 19410 18630 19430
rect 18660 19890 18740 19910
rect 18660 19430 18680 19890
rect 18720 19430 18740 19890
rect 18660 19410 18740 19430
rect 18770 19890 18850 19910
rect 18770 19430 18790 19890
rect 18830 19430 18850 19890
rect 18770 19410 18850 19430
rect 18880 19890 18960 19910
rect 18880 19430 18900 19890
rect 18940 19430 18960 19890
rect 18880 19410 18960 19430
rect 18990 19890 19070 19910
rect 18990 19430 19010 19890
rect 19050 19430 19070 19890
rect 18990 19410 19070 19430
rect 19100 19890 19180 19910
rect 19100 19430 19120 19890
rect 19160 19430 19180 19890
rect 19100 19410 19180 19430
rect 19210 19890 19290 19910
rect 19210 19430 19230 19890
rect 19270 19430 19290 19890
rect 19210 19410 19290 19430
rect 19320 19890 19400 19910
rect 19320 19430 19340 19890
rect 19380 19430 19400 19890
rect 19320 19410 19400 19430
rect 19430 19890 19510 19910
rect 19430 19430 19450 19890
rect 19490 19430 19510 19890
rect 19430 19410 19510 19430
rect 19540 19890 19620 19910
rect 19540 19430 19560 19890
rect 19600 19430 19620 19890
rect 19540 19410 19620 19430
rect 19650 19890 19730 19910
rect 19650 19430 19670 19890
rect 19710 19430 19730 19890
rect 19650 19410 19730 19430
rect 19760 19890 19840 19910
rect 19760 19430 19780 19890
rect 19820 19430 19840 19890
rect 19760 19410 19840 19430
rect 19870 19890 19950 19910
rect 19870 19430 19890 19890
rect 19930 19430 19950 19890
rect 19870 19410 19950 19430
rect 19980 19890 20060 19910
rect 19980 19430 20000 19890
rect 20040 19430 20060 19890
rect 19980 19410 20060 19430
rect 20090 19890 20170 19910
rect 20090 19430 20110 19890
rect 20150 19430 20170 19890
rect 20090 19410 20170 19430
rect 20200 19890 20280 19910
rect 20200 19430 20220 19890
rect 20260 19430 20280 19890
rect 20200 19410 20280 19430
rect 20310 19890 20390 19910
rect 20310 19430 20330 19890
rect 20370 19430 20390 19890
rect 20310 19410 20390 19430
rect 20420 19890 20500 19910
rect 20420 19430 20440 19890
rect 20480 19430 20500 19890
rect 20420 19410 20500 19430
rect 20530 19890 20600 19910
rect 20530 19430 20550 19890
rect 20590 19430 20600 19890
rect 20530 19410 20600 19430
rect 9760 14890 9830 14910
rect 9760 14430 9770 14890
rect 9810 14430 9830 14890
rect 9760 14410 9830 14430
rect 9860 14890 9940 14910
rect 9860 14430 9880 14890
rect 9920 14430 9940 14890
rect 9860 14410 9940 14430
rect 9970 14890 10040 14910
rect 9970 14430 9990 14890
rect 10030 14430 10040 14890
rect 9970 14410 10040 14430
rect 10300 14410 10370 14910
rect 10400 14890 10480 14910
rect 10400 14430 10420 14890
rect 10460 14430 10480 14890
rect 10400 14410 10480 14430
rect 10510 14890 10630 14910
rect 10510 14430 10550 14890
rect 10590 14430 10630 14890
rect 10510 14410 10630 14430
rect 10660 14890 10740 14910
rect 10660 14430 10680 14890
rect 10720 14430 10740 14890
rect 10660 14410 10740 14430
rect 10770 14410 10840 14910
rect 10900 14890 10970 14910
rect 10900 14430 10910 14890
rect 10950 14430 10970 14890
rect 10900 14410 10970 14430
rect 11000 14890 11080 14910
rect 11000 14430 11020 14890
rect 11060 14430 11080 14890
rect 11000 14410 11080 14430
rect 11110 14890 11180 14910
rect 11110 14430 11130 14890
rect 11170 14430 11180 14890
rect 11110 14410 11180 14430
rect 11290 14410 11360 14910
rect 11390 14890 11470 14910
rect 11390 14430 11410 14890
rect 11450 14430 11470 14890
rect 11390 14410 11470 14430
rect 11500 14890 11620 14910
rect 11500 14430 11540 14890
rect 11580 14430 11620 14890
rect 11500 14410 11620 14430
rect 11650 14890 11730 14910
rect 11650 14430 11670 14890
rect 11710 14430 11730 14890
rect 11650 14410 11730 14430
rect 11760 14410 11830 14910
rect 11890 14890 11960 14910
rect 11890 14430 11900 14890
rect 11940 14430 11960 14890
rect 11890 14410 11960 14430
rect 11990 14890 12070 14910
rect 11990 14430 12010 14890
rect 12050 14430 12070 14890
rect 11990 14410 12070 14430
rect 12100 14890 12170 14910
rect 12100 14430 12120 14890
rect 12160 14430 12170 14890
rect 12100 14410 12170 14430
rect 12290 14410 12360 14910
rect 12390 14890 12470 14910
rect 12390 14430 12410 14890
rect 12450 14430 12470 14890
rect 12390 14410 12470 14430
rect 12500 14890 12620 14910
rect 12500 14430 12540 14890
rect 12580 14430 12620 14890
rect 12500 14410 12620 14430
rect 12650 14890 12730 14910
rect 12650 14430 12670 14890
rect 12710 14430 12730 14890
rect 12650 14410 12730 14430
rect 12760 14410 12830 14910
rect 12890 14890 12960 14910
rect 12890 14430 12900 14890
rect 12940 14430 12960 14890
rect 12890 14410 12960 14430
rect 12990 14890 13070 14910
rect 12990 14430 13010 14890
rect 13050 14430 13070 14890
rect 12990 14410 13070 14430
rect 13100 14890 13170 14910
rect 13100 14430 13120 14890
rect 13160 14430 13170 14890
rect 13100 14410 13170 14430
rect 13240 14890 13310 14910
rect 13240 14430 13250 14890
rect 13290 14430 13310 14890
rect 13240 14410 13310 14430
rect 13340 14890 13410 14910
rect 13340 14430 13360 14890
rect 13400 14430 13410 14890
rect 13340 14410 13410 14430
rect 13470 14890 13540 14910
rect 13470 14430 13480 14890
rect 13520 14430 13540 14890
rect 13470 14410 13540 14430
rect 13570 14890 13650 14910
rect 13570 14430 13590 14890
rect 13630 14430 13650 14890
rect 13570 14410 13650 14430
rect 13680 14890 13750 14910
rect 13680 14430 13700 14890
rect 13740 14430 13750 14890
rect 13680 14410 13750 14430
rect 13810 14890 13880 14910
rect 13810 14430 13820 14890
rect 13860 14430 13880 14890
rect 13810 14410 13880 14430
rect 13910 14890 13990 14910
rect 13910 14430 13930 14890
rect 13970 14430 13990 14890
rect 13910 14410 13990 14430
rect 14020 14890 14100 14910
rect 14020 14430 14040 14890
rect 14080 14430 14100 14890
rect 14020 14410 14100 14430
rect 14130 14890 14210 14910
rect 14130 14430 14150 14890
rect 14190 14430 14210 14890
rect 14130 14410 14210 14430
rect 14240 14890 14310 14910
rect 14240 14430 14260 14890
rect 14300 14430 14310 14890
rect 14240 14410 14310 14430
rect 14370 14890 14440 14910
rect 14370 14430 14380 14890
rect 14420 14430 14440 14890
rect 14370 14410 14440 14430
rect 14470 14890 14550 14910
rect 14470 14430 14490 14890
rect 14530 14430 14550 14890
rect 14470 14410 14550 14430
rect 14580 14890 14660 14910
rect 14580 14430 14600 14890
rect 14640 14430 14660 14890
rect 14580 14410 14660 14430
rect 14690 14890 14770 14910
rect 14690 14430 14710 14890
rect 14750 14430 14770 14890
rect 14690 14410 14770 14430
rect 14800 14890 14880 14910
rect 14800 14430 14820 14890
rect 14860 14430 14880 14890
rect 14800 14410 14880 14430
rect 14910 14890 14990 14910
rect 14910 14430 14930 14890
rect 14970 14430 14990 14890
rect 14910 14410 14990 14430
rect 15020 14890 15100 14910
rect 15020 14430 15040 14890
rect 15080 14430 15100 14890
rect 15020 14410 15100 14430
rect 15130 14890 15210 14910
rect 15130 14430 15150 14890
rect 15190 14430 15210 14890
rect 15130 14410 15210 14430
rect 15240 14890 15310 14910
rect 15240 14430 15260 14890
rect 15300 14430 15310 14890
rect 15240 14410 15310 14430
rect 15430 14890 15500 14910
rect 15430 14430 15440 14890
rect 15480 14430 15500 14890
rect 15430 14410 15500 14430
rect 15530 14890 15610 14910
rect 15530 14430 15550 14890
rect 15590 14430 15610 14890
rect 15530 14410 15610 14430
rect 15640 14890 15720 14910
rect 15640 14430 15660 14890
rect 15700 14430 15720 14890
rect 15640 14410 15720 14430
rect 15750 14890 15830 14910
rect 15750 14430 15770 14890
rect 15810 14430 15830 14890
rect 15750 14410 15830 14430
rect 15860 14890 15940 14910
rect 15860 14430 15880 14890
rect 15920 14430 15940 14890
rect 15860 14410 15940 14430
rect 15970 14890 16050 14910
rect 15970 14430 15990 14890
rect 16030 14430 16050 14890
rect 15970 14410 16050 14430
rect 16080 14890 16160 14910
rect 16080 14430 16100 14890
rect 16140 14430 16160 14890
rect 16080 14410 16160 14430
rect 16190 14890 16270 14910
rect 16190 14430 16210 14890
rect 16250 14430 16270 14890
rect 16190 14410 16270 14430
rect 16300 14890 16380 14910
rect 16300 14430 16320 14890
rect 16360 14430 16380 14890
rect 16300 14410 16380 14430
rect 16410 14890 16490 14910
rect 16410 14430 16430 14890
rect 16470 14430 16490 14890
rect 16410 14410 16490 14430
rect 16520 14890 16600 14910
rect 16520 14430 16540 14890
rect 16580 14430 16600 14890
rect 16520 14410 16600 14430
rect 16630 14890 16710 14910
rect 16630 14430 16650 14890
rect 16690 14430 16710 14890
rect 16630 14410 16710 14430
rect 16740 14890 16820 14910
rect 16740 14430 16760 14890
rect 16800 14430 16820 14890
rect 16740 14410 16820 14430
rect 16850 14890 16930 14910
rect 16850 14430 16870 14890
rect 16910 14430 16930 14890
rect 16850 14410 16930 14430
rect 16960 14890 17040 14910
rect 16960 14430 16980 14890
rect 17020 14430 17040 14890
rect 16960 14410 17040 14430
rect 17070 14890 17150 14910
rect 17070 14430 17090 14890
rect 17130 14430 17150 14890
rect 17070 14410 17150 14430
rect 17180 14890 17250 14910
rect 17180 14430 17200 14890
rect 17240 14430 17250 14890
rect 17180 14410 17250 14430
rect 17380 14890 17450 14910
rect 17380 14430 17390 14890
rect 17430 14430 17450 14890
rect 17380 14410 17450 14430
rect 17480 14890 17560 14910
rect 17480 14430 17500 14890
rect 17540 14430 17560 14890
rect 17480 14410 17560 14430
rect 17590 14890 17670 14910
rect 17590 14430 17610 14890
rect 17650 14430 17670 14890
rect 17590 14410 17670 14430
rect 17700 14890 17780 14910
rect 17700 14430 17720 14890
rect 17760 14430 17780 14890
rect 17700 14410 17780 14430
rect 17810 14890 17890 14910
rect 17810 14430 17830 14890
rect 17870 14430 17890 14890
rect 17810 14410 17890 14430
rect 17920 14890 18000 14910
rect 17920 14430 17940 14890
rect 17980 14430 18000 14890
rect 17920 14410 18000 14430
rect 18030 14890 18110 14910
rect 18030 14430 18050 14890
rect 18090 14430 18110 14890
rect 18030 14410 18110 14430
rect 18140 14890 18220 14910
rect 18140 14430 18160 14890
rect 18200 14430 18220 14890
rect 18140 14410 18220 14430
rect 18250 14890 18330 14910
rect 18250 14430 18270 14890
rect 18310 14430 18330 14890
rect 18250 14410 18330 14430
rect 18360 14890 18440 14910
rect 18360 14430 18380 14890
rect 18420 14430 18440 14890
rect 18360 14410 18440 14430
rect 18470 14890 18550 14910
rect 18470 14430 18490 14890
rect 18530 14430 18550 14890
rect 18470 14410 18550 14430
rect 18580 14890 18660 14910
rect 18580 14430 18600 14890
rect 18640 14430 18660 14890
rect 18580 14410 18660 14430
rect 18690 14890 18770 14910
rect 18690 14430 18710 14890
rect 18750 14430 18770 14890
rect 18690 14410 18770 14430
rect 18800 14890 18880 14910
rect 18800 14430 18820 14890
rect 18860 14430 18880 14890
rect 18800 14410 18880 14430
rect 18910 14890 18990 14910
rect 18910 14430 18930 14890
rect 18970 14430 18990 14890
rect 18910 14410 18990 14430
rect 19020 14890 19100 14910
rect 19020 14430 19040 14890
rect 19080 14430 19100 14890
rect 19020 14410 19100 14430
rect 19130 14890 19210 14910
rect 19130 14430 19150 14890
rect 19190 14430 19210 14890
rect 19130 14410 19210 14430
rect 19240 14890 19320 14910
rect 19240 14430 19260 14890
rect 19300 14430 19320 14890
rect 19240 14410 19320 14430
rect 19350 14890 19430 14910
rect 19350 14430 19370 14890
rect 19410 14430 19430 14890
rect 19350 14410 19430 14430
rect 19460 14890 19540 14910
rect 19460 14430 19480 14890
rect 19520 14430 19540 14890
rect 19460 14410 19540 14430
rect 19570 14890 19650 14910
rect 19570 14430 19590 14890
rect 19630 14430 19650 14890
rect 19570 14410 19650 14430
rect 19680 14890 19760 14910
rect 19680 14430 19700 14890
rect 19740 14430 19760 14890
rect 19680 14410 19760 14430
rect 19790 14890 19870 14910
rect 19790 14430 19810 14890
rect 19850 14430 19870 14890
rect 19790 14410 19870 14430
rect 19900 14890 19980 14910
rect 19900 14430 19920 14890
rect 19960 14430 19980 14890
rect 19900 14410 19980 14430
rect 20010 14890 20090 14910
rect 20010 14430 20030 14890
rect 20070 14430 20090 14890
rect 20010 14410 20090 14430
rect 20120 14890 20200 14910
rect 20120 14430 20140 14890
rect 20180 14430 20200 14890
rect 20120 14410 20200 14430
rect 20230 14890 20310 14910
rect 20230 14430 20250 14890
rect 20290 14430 20310 14890
rect 20230 14410 20310 14430
rect 20340 14890 20420 14910
rect 20340 14430 20360 14890
rect 20400 14430 20420 14890
rect 20340 14410 20420 14430
rect 20450 14890 20530 14910
rect 20450 14430 20470 14890
rect 20510 14430 20530 14890
rect 20450 14410 20530 14430
rect 20560 14890 20640 14910
rect 20560 14430 20580 14890
rect 20620 14430 20640 14890
rect 20560 14410 20640 14430
rect 20670 14890 20750 14910
rect 20670 14430 20690 14890
rect 20730 14430 20750 14890
rect 20670 14410 20750 14430
rect 20780 14890 20860 14910
rect 20780 14430 20800 14890
rect 20840 14430 20860 14890
rect 20780 14410 20860 14430
rect 20890 14890 20960 14910
rect 20890 14430 20910 14890
rect 20950 14430 20960 14890
rect 20890 14410 20960 14430
rect 7280 13240 7350 13260
rect 7280 12780 7290 13240
rect 7330 12780 7350 13240
rect 7280 12760 7350 12780
rect 7380 13240 7460 13260
rect 7380 12780 7400 13240
rect 7440 12780 7460 13240
rect 7380 12760 7460 12780
rect 7490 13240 7560 13260
rect 7490 12780 7510 13240
rect 7550 12780 7560 13240
rect 7490 12760 7560 12780
rect 7800 12760 7870 13260
rect 7900 13240 7980 13260
rect 7900 12780 7920 13240
rect 7960 12780 7980 13240
rect 7900 12760 7980 12780
rect 8010 13240 8130 13260
rect 8010 12780 8050 13240
rect 8090 12780 8130 13240
rect 8010 12760 8130 12780
rect 8160 13240 8240 13260
rect 8160 12780 8180 13240
rect 8220 12780 8240 13240
rect 8160 12760 8240 12780
rect 8270 12760 8340 13260
rect 8550 13240 8620 13260
rect 8550 12780 8560 13240
rect 8600 12780 8620 13240
rect 8550 12760 8620 12780
rect 8650 13240 8770 13260
rect 8650 12780 8690 13240
rect 8730 12780 8770 13240
rect 8650 12760 8770 12780
rect 8800 13240 8870 13260
rect 8800 12780 8820 13240
rect 8860 12780 8870 13240
rect 8800 12760 8870 12780
rect 8930 13240 9000 13260
rect 8930 12780 8940 13240
rect 8980 12780 9000 13240
rect 8930 12760 9000 12780
rect 9030 13240 9100 13260
rect 9030 12780 9050 13240
rect 9090 12780 9100 13240
rect 9030 12760 9100 12780
rect 9190 13240 9260 13260
rect 9190 12780 9200 13240
rect 9240 12780 9260 13240
rect 9190 12760 9260 12780
rect 9290 13240 9360 13260
rect 9290 12780 9310 13240
rect 9350 12780 9360 13240
rect 9290 12760 9360 12780
rect 9440 13240 9510 13260
rect 9440 12780 9450 13240
rect 9490 12780 9510 13240
rect 9440 12760 9510 12780
rect 9540 13240 9610 13260
rect 9540 12780 9560 13240
rect 9600 12780 9610 13240
rect 9540 12760 9610 12780
rect 9860 13240 9930 13260
rect 9860 12780 9870 13240
rect 9910 12780 9930 13240
rect 9860 12760 9930 12780
rect 9960 13240 10040 13260
rect 9960 12780 9980 13240
rect 10020 12780 10040 13240
rect 9960 12760 10040 12780
rect 10070 13240 10140 13260
rect 10070 12780 10090 13240
rect 10130 12780 10140 13240
rect 10070 12760 10140 12780
rect 10400 12760 10470 13260
rect 10500 13240 10580 13260
rect 10500 12780 10520 13240
rect 10560 12780 10580 13240
rect 10500 12760 10580 12780
rect 10610 13240 10730 13260
rect 10610 12780 10650 13240
rect 10690 12780 10730 13240
rect 10610 12760 10730 12780
rect 10760 13240 10840 13260
rect 10760 12780 10780 13240
rect 10820 12780 10840 13240
rect 10760 12760 10840 12780
rect 10870 12760 10940 13260
rect 11000 13240 11070 13260
rect 11000 12780 11010 13240
rect 11050 12780 11070 13240
rect 11000 12760 11070 12780
rect 11100 13240 11180 13260
rect 11100 12780 11120 13240
rect 11160 12780 11180 13240
rect 11100 12760 11180 12780
rect 11210 13240 11280 13260
rect 11210 12780 11230 13240
rect 11270 12780 11280 13240
rect 11210 12760 11280 12780
rect 11390 12760 11460 13260
rect 11490 13240 11570 13260
rect 11490 12780 11510 13240
rect 11550 12780 11570 13240
rect 11490 12760 11570 12780
rect 11600 13240 11720 13260
rect 11600 12780 11640 13240
rect 11680 12780 11720 13240
rect 11600 12760 11720 12780
rect 11750 13240 11830 13260
rect 11750 12780 11770 13240
rect 11810 12780 11830 13240
rect 11750 12760 11830 12780
rect 11860 12760 11930 13260
rect 11990 13240 12060 13260
rect 11990 12780 12000 13240
rect 12040 12780 12060 13240
rect 11990 12760 12060 12780
rect 12090 13240 12170 13260
rect 12090 12780 12110 13240
rect 12150 12780 12170 13240
rect 12090 12760 12170 12780
rect 12200 13240 12270 13260
rect 12200 12780 12220 13240
rect 12260 12780 12270 13240
rect 12200 12760 12270 12780
rect 12390 12760 12460 13260
rect 12490 13240 12570 13260
rect 12490 12780 12510 13240
rect 12550 12780 12570 13240
rect 12490 12760 12570 12780
rect 12600 13240 12720 13260
rect 12600 12780 12640 13240
rect 12680 12780 12720 13240
rect 12600 12760 12720 12780
rect 12750 13240 12830 13260
rect 12750 12780 12770 13240
rect 12810 12780 12830 13240
rect 12750 12760 12830 12780
rect 12860 12760 12930 13260
rect 12990 13240 13060 13260
rect 12990 12780 13000 13240
rect 13040 12780 13060 13240
rect 12990 12760 13060 12780
rect 13090 13240 13170 13260
rect 13090 12780 13110 13240
rect 13150 12780 13170 13240
rect 13090 12760 13170 12780
rect 13200 13240 13270 13260
rect 13200 12780 13220 13240
rect 13260 12780 13270 13240
rect 13200 12760 13270 12780
rect 13340 13240 13410 13260
rect 13340 12780 13350 13240
rect 13390 12780 13410 13240
rect 13340 12760 13410 12780
rect 13440 13240 13510 13260
rect 13440 12780 13460 13240
rect 13500 12780 13510 13240
rect 13440 12760 13510 12780
rect 13570 13240 13640 13260
rect 13570 12780 13580 13240
rect 13620 12780 13640 13240
rect 13570 12760 13640 12780
rect 13670 13240 13750 13260
rect 13670 12780 13690 13240
rect 13730 12780 13750 13240
rect 13670 12760 13750 12780
rect 13780 13240 13850 13260
rect 13780 12780 13800 13240
rect 13840 12780 13850 13240
rect 13780 12760 13850 12780
rect 13910 13240 13980 13260
rect 13910 12780 13920 13240
rect 13960 12780 13980 13240
rect 13910 12760 13980 12780
rect 14010 13240 14090 13260
rect 14010 12780 14030 13240
rect 14070 12780 14090 13240
rect 14010 12760 14090 12780
rect 14120 13240 14200 13260
rect 14120 12780 14140 13240
rect 14180 12780 14200 13240
rect 14120 12760 14200 12780
rect 14230 13240 14310 13260
rect 14230 12780 14250 13240
rect 14290 12780 14310 13240
rect 14230 12760 14310 12780
rect 14340 13240 14410 13260
rect 14340 12780 14360 13240
rect 14400 12780 14410 13240
rect 14340 12760 14410 12780
rect 14470 13240 14540 13260
rect 14470 12780 14480 13240
rect 14520 12780 14540 13240
rect 14470 12760 14540 12780
rect 14570 13240 14650 13260
rect 14570 12780 14590 13240
rect 14630 12780 14650 13240
rect 14570 12760 14650 12780
rect 14680 13240 14760 13260
rect 14680 12780 14700 13240
rect 14740 12780 14760 13240
rect 14680 12760 14760 12780
rect 14790 13240 14870 13260
rect 14790 12780 14810 13240
rect 14850 12780 14870 13240
rect 14790 12760 14870 12780
rect 14900 13240 14980 13260
rect 14900 12780 14920 13240
rect 14960 12780 14980 13240
rect 14900 12760 14980 12780
rect 15010 13240 15090 13260
rect 15010 12780 15030 13240
rect 15070 12780 15090 13240
rect 15010 12760 15090 12780
rect 15120 13240 15200 13260
rect 15120 12780 15140 13240
rect 15180 12780 15200 13240
rect 15120 12760 15200 12780
rect 15230 13240 15310 13260
rect 15230 12780 15250 13240
rect 15290 12780 15310 13240
rect 15230 12760 15310 12780
rect 15340 13240 15410 13260
rect 15340 12780 15360 13240
rect 15400 12780 15410 13240
rect 15340 12760 15410 12780
rect 15530 13240 15600 13260
rect 15530 12780 15540 13240
rect 15580 12780 15600 13240
rect 15530 12760 15600 12780
rect 15630 13240 15710 13260
rect 15630 12780 15650 13240
rect 15690 12780 15710 13240
rect 15630 12760 15710 12780
rect 15740 13240 15820 13260
rect 15740 12780 15760 13240
rect 15800 12780 15820 13240
rect 15740 12760 15820 12780
rect 15850 13240 15930 13260
rect 15850 12780 15870 13240
rect 15910 12780 15930 13240
rect 15850 12760 15930 12780
rect 15960 13240 16040 13260
rect 15960 12780 15980 13240
rect 16020 12780 16040 13240
rect 15960 12760 16040 12780
rect 16070 13240 16150 13260
rect 16070 12780 16090 13240
rect 16130 12780 16150 13240
rect 16070 12760 16150 12780
rect 16180 13240 16260 13260
rect 16180 12780 16200 13240
rect 16240 12780 16260 13240
rect 16180 12760 16260 12780
rect 16290 13240 16370 13260
rect 16290 12780 16310 13240
rect 16350 12780 16370 13240
rect 16290 12760 16370 12780
rect 16400 13240 16480 13260
rect 16400 12780 16420 13240
rect 16460 12780 16480 13240
rect 16400 12760 16480 12780
rect 16510 13240 16590 13260
rect 16510 12780 16530 13240
rect 16570 12780 16590 13240
rect 16510 12760 16590 12780
rect 16620 13240 16700 13260
rect 16620 12780 16640 13240
rect 16680 12780 16700 13240
rect 16620 12760 16700 12780
rect 16730 13240 16810 13260
rect 16730 12780 16750 13240
rect 16790 12780 16810 13240
rect 16730 12760 16810 12780
rect 16840 13240 16920 13260
rect 16840 12780 16860 13240
rect 16900 12780 16920 13240
rect 16840 12760 16920 12780
rect 16950 13240 17030 13260
rect 16950 12780 16970 13240
rect 17010 12780 17030 13240
rect 16950 12760 17030 12780
rect 17060 13240 17140 13260
rect 17060 12780 17080 13240
rect 17120 12780 17140 13240
rect 17060 12760 17140 12780
rect 17170 13240 17250 13260
rect 17170 12780 17190 13240
rect 17230 12780 17250 13240
rect 17170 12760 17250 12780
rect 17280 13240 17350 13260
rect 17280 12780 17300 13240
rect 17340 12780 17350 13240
rect 17280 12760 17350 12780
rect 17480 13240 17550 13260
rect 17480 12780 17490 13240
rect 17530 12780 17550 13240
rect 17480 12760 17550 12780
rect 17580 13240 17660 13260
rect 17580 12780 17600 13240
rect 17640 12780 17660 13240
rect 17580 12760 17660 12780
rect 17690 13240 17770 13260
rect 17690 12780 17710 13240
rect 17750 12780 17770 13240
rect 17690 12760 17770 12780
rect 17800 13240 17880 13260
rect 17800 12780 17820 13240
rect 17860 12780 17880 13240
rect 17800 12760 17880 12780
rect 17910 13240 17990 13260
rect 17910 12780 17930 13240
rect 17970 12780 17990 13240
rect 17910 12760 17990 12780
rect 18020 13240 18100 13260
rect 18020 12780 18040 13240
rect 18080 12780 18100 13240
rect 18020 12760 18100 12780
rect 18130 13240 18210 13260
rect 18130 12780 18150 13240
rect 18190 12780 18210 13240
rect 18130 12760 18210 12780
rect 18240 13240 18320 13260
rect 18240 12780 18260 13240
rect 18300 12780 18320 13240
rect 18240 12760 18320 12780
rect 18350 13240 18430 13260
rect 18350 12780 18370 13240
rect 18410 12780 18430 13240
rect 18350 12760 18430 12780
rect 18460 13240 18540 13260
rect 18460 12780 18480 13240
rect 18520 12780 18540 13240
rect 18460 12760 18540 12780
rect 18570 13240 18650 13260
rect 18570 12780 18590 13240
rect 18630 12780 18650 13240
rect 18570 12760 18650 12780
rect 18680 13240 18760 13260
rect 18680 12780 18700 13240
rect 18740 12780 18760 13240
rect 18680 12760 18760 12780
rect 18790 13240 18870 13260
rect 18790 12780 18810 13240
rect 18850 12780 18870 13240
rect 18790 12760 18870 12780
rect 18900 13240 18980 13260
rect 18900 12780 18920 13240
rect 18960 12780 18980 13240
rect 18900 12760 18980 12780
rect 19010 13240 19090 13260
rect 19010 12780 19030 13240
rect 19070 12780 19090 13240
rect 19010 12760 19090 12780
rect 19120 13240 19200 13260
rect 19120 12780 19140 13240
rect 19180 12780 19200 13240
rect 19120 12760 19200 12780
rect 19230 13240 19310 13260
rect 19230 12780 19250 13240
rect 19290 12780 19310 13240
rect 19230 12760 19310 12780
rect 19340 13240 19420 13260
rect 19340 12780 19360 13240
rect 19400 12780 19420 13240
rect 19340 12760 19420 12780
rect 19450 13240 19530 13260
rect 19450 12780 19470 13240
rect 19510 12780 19530 13240
rect 19450 12760 19530 12780
rect 19560 13240 19640 13260
rect 19560 12780 19580 13240
rect 19620 12780 19640 13240
rect 19560 12760 19640 12780
rect 19670 13240 19750 13260
rect 19670 12780 19690 13240
rect 19730 12780 19750 13240
rect 19670 12760 19750 12780
rect 19780 13240 19860 13260
rect 19780 12780 19800 13240
rect 19840 12780 19860 13240
rect 19780 12760 19860 12780
rect 19890 13240 19970 13260
rect 19890 12780 19910 13240
rect 19950 12780 19970 13240
rect 19890 12760 19970 12780
rect 20000 13240 20080 13260
rect 20000 12780 20020 13240
rect 20060 12780 20080 13240
rect 20000 12760 20080 12780
rect 20110 13240 20190 13260
rect 20110 12780 20130 13240
rect 20170 12780 20190 13240
rect 20110 12760 20190 12780
rect 20220 13240 20300 13260
rect 20220 12780 20240 13240
rect 20280 12780 20300 13240
rect 20220 12760 20300 12780
rect 20330 13240 20410 13260
rect 20330 12780 20350 13240
rect 20390 12780 20410 13240
rect 20330 12760 20410 12780
rect 20440 13240 20520 13260
rect 20440 12780 20460 13240
rect 20500 12780 20520 13240
rect 20440 12760 20520 12780
rect 20550 13240 20630 13260
rect 20550 12780 20570 13240
rect 20610 12780 20630 13240
rect 20550 12760 20630 12780
rect 20660 13240 20740 13260
rect 20660 12780 20680 13240
rect 20720 12780 20740 13240
rect 20660 12760 20740 12780
rect 20770 13240 20850 13260
rect 20770 12780 20790 13240
rect 20830 12780 20850 13240
rect 20770 12760 20850 12780
rect 20880 13240 20960 13260
rect 20880 12780 20900 13240
rect 20940 12780 20960 13240
rect 20880 12760 20960 12780
rect 20990 13240 21060 13260
rect 20990 12780 21010 13240
rect 21050 12780 21060 13240
rect 20990 12760 21060 12780
rect 7280 10270 7350 10290
rect 7280 9810 7290 10270
rect 7330 9810 7350 10270
rect 7280 9790 7350 9810
rect 7380 10270 7460 10290
rect 7380 9810 7400 10270
rect 7440 9810 7460 10270
rect 7380 9790 7460 9810
rect 7490 10270 7560 10290
rect 7490 9810 7510 10270
rect 7550 9810 7560 10270
rect 7490 9790 7560 9810
rect 7850 9720 7920 10720
rect 7950 10700 8030 10720
rect 7950 9740 7970 10700
rect 8010 9740 8030 10700
rect 7950 9720 8030 9740
rect 8060 9720 8180 10720
rect 8210 10700 8290 10720
rect 8210 9740 8230 10700
rect 8270 9740 8290 10700
rect 8210 9720 8290 9740
rect 8320 9720 8390 10720
rect 8640 10280 8710 10300
rect 8640 9820 8650 10280
rect 8690 9820 8710 10280
rect 8640 9800 8710 9820
rect 8740 10280 8860 10300
rect 8740 9820 8780 10280
rect 8820 9820 8860 10280
rect 8740 9800 8860 9820
rect 8890 10280 8960 10300
rect 8890 9820 8910 10280
rect 8950 9820 8960 10280
rect 8890 9800 8960 9820
rect 9020 10280 9090 10300
rect 9020 9820 9030 10280
rect 9070 9820 9090 10280
rect 9020 9800 9090 9820
rect 9120 10280 9190 10300
rect 9120 9820 9140 10280
rect 9180 9820 9190 10280
rect 9120 9800 9190 9820
rect 9280 10280 9350 10300
rect 9280 9820 9290 10280
rect 9330 9820 9350 10280
rect 9280 9800 9350 9820
rect 9380 10280 9450 10300
rect 9380 9820 9400 10280
rect 9440 9820 9450 10280
rect 9380 9800 9450 9820
rect 9530 10280 9600 10300
rect 9530 9820 9540 10280
rect 9580 9820 9600 10280
rect 9530 9800 9600 9820
rect 9630 10280 9700 10300
rect 9630 9820 9650 10280
rect 9690 9820 9700 10280
rect 9630 9800 9700 9820
rect 9860 10270 9930 10290
rect 9860 9810 9870 10270
rect 9910 9810 9930 10270
rect 9860 9790 9930 9810
rect 9960 10270 10040 10290
rect 9960 9810 9980 10270
rect 10020 9810 10040 10270
rect 9960 9790 10040 9810
rect 10070 10270 10140 10290
rect 10070 9810 10090 10270
rect 10130 9810 10140 10270
rect 10070 9790 10140 9810
rect 10400 9790 10470 10290
rect 10500 10270 10580 10290
rect 10500 9810 10520 10270
rect 10560 9810 10580 10270
rect 10500 9790 10580 9810
rect 10610 10270 10730 10290
rect 10610 9810 10650 10270
rect 10690 9810 10730 10270
rect 10610 9790 10730 9810
rect 10760 10270 10840 10290
rect 10760 9810 10780 10270
rect 10820 9810 10840 10270
rect 10760 9790 10840 9810
rect 10870 9790 10940 10290
rect 11000 10270 11070 10290
rect 11000 9810 11010 10270
rect 11050 9810 11070 10270
rect 11000 9790 11070 9810
rect 11100 10270 11180 10290
rect 11100 9810 11120 10270
rect 11160 9810 11180 10270
rect 11100 9790 11180 9810
rect 11210 10270 11280 10290
rect 11210 9810 11230 10270
rect 11270 9810 11280 10270
rect 11210 9790 11280 9810
rect 11390 9790 11460 10290
rect 11490 10270 11570 10290
rect 11490 9810 11510 10270
rect 11550 9810 11570 10270
rect 11490 9790 11570 9810
rect 11600 10270 11720 10290
rect 11600 9810 11640 10270
rect 11680 9810 11720 10270
rect 11600 9790 11720 9810
rect 11750 10270 11830 10290
rect 11750 9810 11770 10270
rect 11810 9810 11830 10270
rect 11750 9790 11830 9810
rect 11860 9790 11930 10290
rect 11990 10270 12060 10290
rect 11990 9810 12000 10270
rect 12040 9810 12060 10270
rect 11990 9790 12060 9810
rect 12090 10270 12170 10290
rect 12090 9810 12110 10270
rect 12150 9810 12170 10270
rect 12090 9790 12170 9810
rect 12200 10270 12270 10290
rect 12200 9810 12220 10270
rect 12260 9810 12270 10270
rect 12200 9790 12270 9810
rect 12390 9790 12460 10290
rect 12490 10270 12570 10290
rect 12490 9810 12510 10270
rect 12550 9810 12570 10270
rect 12490 9790 12570 9810
rect 12600 10270 12720 10290
rect 12600 9810 12640 10270
rect 12680 9810 12720 10270
rect 12600 9790 12720 9810
rect 12750 10270 12830 10290
rect 12750 9810 12770 10270
rect 12810 9810 12830 10270
rect 12750 9790 12830 9810
rect 12860 9790 12930 10290
rect 12990 10270 13060 10290
rect 12990 9810 13000 10270
rect 13040 9810 13060 10270
rect 12990 9790 13060 9810
rect 13090 10270 13170 10290
rect 13090 9810 13110 10270
rect 13150 9810 13170 10270
rect 13090 9790 13170 9810
rect 13200 10270 13270 10290
rect 13200 9810 13220 10270
rect 13260 9810 13270 10270
rect 13200 9790 13270 9810
rect 13330 10270 13400 10290
rect 13330 9810 13340 10270
rect 13380 9810 13400 10270
rect 13330 9790 13400 9810
rect 13430 10270 13500 10290
rect 13430 9810 13450 10270
rect 13490 9810 13500 10270
rect 13430 9790 13500 9810
rect 13560 10270 13630 10290
rect 13560 9810 13570 10270
rect 13610 9810 13630 10270
rect 13560 9790 13630 9810
rect 13660 10270 13740 10290
rect 13660 9810 13680 10270
rect 13720 9810 13740 10270
rect 13660 9790 13740 9810
rect 13770 10270 13840 10290
rect 13770 9810 13790 10270
rect 13830 9810 13840 10270
rect 13770 9790 13840 9810
rect 13900 10270 13970 10290
rect 13900 9810 13910 10270
rect 13950 9810 13970 10270
rect 13900 9790 13970 9810
rect 14000 10270 14080 10290
rect 14000 9810 14020 10270
rect 14060 9810 14080 10270
rect 14000 9790 14080 9810
rect 14110 10270 14190 10290
rect 14110 9810 14130 10270
rect 14170 9810 14190 10270
rect 14110 9790 14190 9810
rect 14220 10270 14300 10290
rect 14220 9810 14240 10270
rect 14280 9810 14300 10270
rect 14220 9790 14300 9810
rect 14330 10270 14400 10290
rect 14330 9810 14350 10270
rect 14390 9810 14400 10270
rect 14330 9790 14400 9810
rect 14460 10270 14530 10290
rect 14460 9810 14470 10270
rect 14510 9810 14530 10270
rect 14460 9790 14530 9810
rect 14560 10270 14640 10290
rect 14560 9810 14580 10270
rect 14620 9810 14640 10270
rect 14560 9790 14640 9810
rect 14670 10270 14750 10290
rect 14670 9810 14690 10270
rect 14730 9810 14750 10270
rect 14670 9790 14750 9810
rect 14780 10270 14860 10290
rect 14780 9810 14800 10270
rect 14840 9810 14860 10270
rect 14780 9790 14860 9810
rect 14890 10270 14970 10290
rect 14890 9810 14910 10270
rect 14950 9810 14970 10270
rect 14890 9790 14970 9810
rect 15000 10270 15080 10290
rect 15000 9810 15020 10270
rect 15060 9810 15080 10270
rect 15000 9790 15080 9810
rect 15110 10270 15190 10290
rect 15110 9810 15130 10270
rect 15170 9810 15190 10270
rect 15110 9790 15190 9810
rect 15220 10270 15300 10290
rect 15220 9810 15240 10270
rect 15280 9810 15300 10270
rect 15220 9790 15300 9810
rect 15330 10270 15400 10290
rect 15330 9810 15350 10270
rect 15390 9810 15400 10270
rect 15330 9790 15400 9810
rect 15520 10270 15590 10290
rect 15520 9810 15530 10270
rect 15570 9810 15590 10270
rect 15520 9790 15590 9810
rect 15620 10270 15700 10290
rect 15620 9810 15640 10270
rect 15680 9810 15700 10270
rect 15620 9790 15700 9810
rect 15730 10270 15810 10290
rect 15730 9810 15750 10270
rect 15790 9810 15810 10270
rect 15730 9790 15810 9810
rect 15840 10270 15920 10290
rect 15840 9810 15860 10270
rect 15900 9810 15920 10270
rect 15840 9790 15920 9810
rect 15950 10270 16030 10290
rect 15950 9810 15970 10270
rect 16010 9810 16030 10270
rect 15950 9790 16030 9810
rect 16060 10270 16140 10290
rect 16060 9810 16080 10270
rect 16120 9810 16140 10270
rect 16060 9790 16140 9810
rect 16170 10270 16250 10290
rect 16170 9810 16190 10270
rect 16230 9810 16250 10270
rect 16170 9790 16250 9810
rect 16280 10270 16360 10290
rect 16280 9810 16300 10270
rect 16340 9810 16360 10270
rect 16280 9790 16360 9810
rect 16390 10270 16470 10290
rect 16390 9810 16410 10270
rect 16450 9810 16470 10270
rect 16390 9790 16470 9810
rect 16500 10270 16580 10290
rect 16500 9810 16520 10270
rect 16560 9810 16580 10270
rect 16500 9790 16580 9810
rect 16610 10270 16690 10290
rect 16610 9810 16630 10270
rect 16670 9810 16690 10270
rect 16610 9790 16690 9810
rect 16720 10270 16800 10290
rect 16720 9810 16740 10270
rect 16780 9810 16800 10270
rect 16720 9790 16800 9810
rect 16830 10270 16910 10290
rect 16830 9810 16850 10270
rect 16890 9810 16910 10270
rect 16830 9790 16910 9810
rect 16940 10270 17020 10290
rect 16940 9810 16960 10270
rect 17000 9810 17020 10270
rect 16940 9790 17020 9810
rect 17050 10270 17130 10290
rect 17050 9810 17070 10270
rect 17110 9810 17130 10270
rect 17050 9790 17130 9810
rect 17160 10270 17240 10290
rect 17160 9810 17180 10270
rect 17220 9810 17240 10270
rect 17160 9790 17240 9810
rect 17270 10270 17340 10290
rect 17270 9810 17290 10270
rect 17330 9810 17340 10270
rect 17270 9790 17340 9810
rect 17470 10270 17540 10290
rect 17470 9810 17480 10270
rect 17520 9810 17540 10270
rect 17470 9790 17540 9810
rect 17570 10270 17650 10290
rect 17570 9810 17590 10270
rect 17630 9810 17650 10270
rect 17570 9790 17650 9810
rect 17680 10270 17760 10290
rect 17680 9810 17700 10270
rect 17740 9810 17760 10270
rect 17680 9790 17760 9810
rect 17790 10270 17870 10290
rect 17790 9810 17810 10270
rect 17850 9810 17870 10270
rect 17790 9790 17870 9810
rect 17900 10270 17980 10290
rect 17900 9810 17920 10270
rect 17960 9810 17980 10270
rect 17900 9790 17980 9810
rect 18010 10270 18090 10290
rect 18010 9810 18030 10270
rect 18070 9810 18090 10270
rect 18010 9790 18090 9810
rect 18120 10270 18200 10290
rect 18120 9810 18140 10270
rect 18180 9810 18200 10270
rect 18120 9790 18200 9810
rect 18230 10270 18310 10290
rect 18230 9810 18250 10270
rect 18290 9810 18310 10270
rect 18230 9790 18310 9810
rect 18340 10270 18420 10290
rect 18340 9810 18360 10270
rect 18400 9810 18420 10270
rect 18340 9790 18420 9810
rect 18450 10270 18530 10290
rect 18450 9810 18470 10270
rect 18510 9810 18530 10270
rect 18450 9790 18530 9810
rect 18560 10270 18640 10290
rect 18560 9810 18580 10270
rect 18620 9810 18640 10270
rect 18560 9790 18640 9810
rect 18670 10270 18750 10290
rect 18670 9810 18690 10270
rect 18730 9810 18750 10270
rect 18670 9790 18750 9810
rect 18780 10270 18860 10290
rect 18780 9810 18800 10270
rect 18840 9810 18860 10270
rect 18780 9790 18860 9810
rect 18890 10270 18970 10290
rect 18890 9810 18910 10270
rect 18950 9810 18970 10270
rect 18890 9790 18970 9810
rect 19000 10270 19080 10290
rect 19000 9810 19020 10270
rect 19060 9810 19080 10270
rect 19000 9790 19080 9810
rect 19110 10270 19190 10290
rect 19110 9810 19130 10270
rect 19170 9810 19190 10270
rect 19110 9790 19190 9810
rect 19220 10270 19300 10290
rect 19220 9810 19240 10270
rect 19280 9810 19300 10270
rect 19220 9790 19300 9810
rect 19330 10270 19410 10290
rect 19330 9810 19350 10270
rect 19390 9810 19410 10270
rect 19330 9790 19410 9810
rect 19440 10270 19520 10290
rect 19440 9810 19460 10270
rect 19500 9810 19520 10270
rect 19440 9790 19520 9810
rect 19550 10270 19630 10290
rect 19550 9810 19570 10270
rect 19610 9810 19630 10270
rect 19550 9790 19630 9810
rect 19660 10270 19740 10290
rect 19660 9810 19680 10270
rect 19720 9810 19740 10270
rect 19660 9790 19740 9810
rect 19770 10270 19850 10290
rect 19770 9810 19790 10270
rect 19830 9810 19850 10270
rect 19770 9790 19850 9810
rect 19880 10270 19960 10290
rect 19880 9810 19900 10270
rect 19940 9810 19960 10270
rect 19880 9790 19960 9810
rect 19990 10270 20070 10290
rect 19990 9810 20010 10270
rect 20050 9810 20070 10270
rect 19990 9790 20070 9810
rect 20100 10270 20180 10290
rect 20100 9810 20120 10270
rect 20160 9810 20180 10270
rect 20100 9790 20180 9810
rect 20210 10270 20290 10290
rect 20210 9810 20230 10270
rect 20270 9810 20290 10270
rect 20210 9790 20290 9810
rect 20320 10270 20400 10290
rect 20320 9810 20340 10270
rect 20380 9810 20400 10270
rect 20320 9790 20400 9810
rect 20430 10270 20510 10290
rect 20430 9810 20450 10270
rect 20490 9810 20510 10270
rect 20430 9790 20510 9810
rect 20540 10270 20620 10290
rect 20540 9810 20560 10270
rect 20600 9810 20620 10270
rect 20540 9790 20620 9810
rect 20650 10270 20730 10290
rect 20650 9810 20670 10270
rect 20710 9810 20730 10270
rect 20650 9790 20730 9810
rect 20760 10270 20840 10290
rect 20760 9810 20780 10270
rect 20820 9810 20840 10270
rect 20760 9790 20840 9810
rect 20870 10270 20950 10290
rect 20870 9810 20890 10270
rect 20930 9810 20950 10270
rect 20870 9790 20950 9810
rect 20980 10270 21050 10290
rect 20980 9810 21000 10270
rect 21040 9810 21050 10270
rect 20980 9790 21050 9810
rect 9900 8240 9970 8260
rect 9900 7080 9910 8240
rect 9950 7080 9970 8240
rect 9900 7060 9970 7080
rect 10000 8240 10080 8260
rect 10000 7080 10020 8240
rect 10060 7080 10080 8240
rect 10000 7060 10080 7080
rect 10110 8240 10190 8260
rect 10110 7080 10130 8240
rect 10170 7080 10190 8240
rect 10110 7060 10190 7080
rect 10220 8240 10300 8260
rect 10220 7080 10240 8240
rect 10280 7080 10300 8240
rect 10220 7060 10300 7080
rect 10330 8240 10410 8260
rect 10330 7080 10350 8240
rect 10390 7080 10410 8240
rect 10330 7060 10410 7080
rect 10440 8240 10520 8260
rect 10440 7080 10460 8240
rect 10500 7080 10520 8240
rect 10440 7060 10520 7080
rect 10550 8240 10630 8260
rect 10550 7080 10570 8240
rect 10610 7080 10630 8240
rect 10550 7060 10630 7080
rect 10660 8240 10740 8260
rect 10660 7080 10680 8240
rect 10720 7080 10740 8240
rect 10660 7060 10740 7080
rect 10770 8240 10850 8260
rect 10770 7080 10790 8240
rect 10830 7080 10850 8240
rect 10770 7060 10850 7080
rect 10880 8240 10960 8260
rect 10880 7080 10900 8240
rect 10940 7080 10960 8240
rect 10880 7060 10960 7080
rect 10990 8240 11070 8260
rect 10990 7080 11010 8240
rect 11050 7080 11070 8240
rect 10990 7060 11070 7080
rect 11100 8240 11180 8260
rect 11100 7080 11120 8240
rect 11160 7080 11180 8240
rect 11100 7060 11180 7080
rect 11210 8240 11290 8260
rect 11210 7080 11230 8240
rect 11270 7080 11290 8240
rect 11210 7060 11290 7080
rect 11320 8240 11400 8260
rect 11320 7080 11340 8240
rect 11380 7080 11400 8240
rect 11320 7060 11400 7080
rect 11430 8240 11510 8260
rect 11430 7080 11450 8240
rect 11490 7080 11510 8240
rect 11430 7060 11510 7080
rect 11540 8240 11620 8260
rect 11540 7080 11560 8240
rect 11600 7080 11620 8240
rect 11540 7060 11620 7080
rect 11650 8240 11730 8260
rect 11650 7080 11670 8240
rect 11710 7080 11730 8240
rect 11650 7060 11730 7080
rect 11760 8240 11840 8260
rect 11760 7080 11780 8240
rect 11820 7080 11840 8240
rect 11760 7060 11840 7080
rect 11870 8240 11950 8260
rect 11870 7080 11890 8240
rect 11930 7080 11950 8240
rect 11870 7060 11950 7080
rect 11980 8240 12060 8260
rect 11980 7080 12000 8240
rect 12040 7080 12060 8240
rect 11980 7060 12060 7080
rect 12090 8240 12170 8260
rect 12090 7080 12110 8240
rect 12150 7080 12170 8240
rect 12090 7060 12170 7080
rect 12200 8240 12280 8260
rect 12200 7080 12220 8240
rect 12260 7080 12280 8240
rect 12200 7060 12280 7080
rect 12310 8240 12390 8260
rect 12310 7080 12330 8240
rect 12370 7080 12390 8240
rect 12310 7060 12390 7080
rect 12420 8240 12500 8260
rect 12420 7080 12440 8240
rect 12480 7080 12500 8240
rect 12420 7060 12500 7080
rect 12530 8240 12610 8260
rect 12530 7080 12550 8240
rect 12590 7080 12610 8240
rect 12530 7060 12610 7080
rect 12640 8240 12720 8260
rect 12640 7080 12660 8240
rect 12700 7080 12720 8240
rect 12640 7060 12720 7080
rect 12750 8240 12830 8260
rect 12750 7080 12770 8240
rect 12810 7080 12830 8240
rect 12750 7060 12830 7080
rect 12860 8240 12940 8260
rect 12860 7080 12880 8240
rect 12920 7080 12940 8240
rect 12860 7060 12940 7080
rect 12970 8240 13050 8260
rect 12970 7080 12990 8240
rect 13030 7080 13050 8240
rect 12970 7060 13050 7080
rect 13080 8240 13160 8260
rect 13080 7080 13100 8240
rect 13140 7080 13160 8240
rect 13080 7060 13160 7080
rect 13190 8240 13260 8260
rect 13190 7080 13210 8240
rect 13250 7080 13260 8240
rect 13190 7060 13260 7080
rect 13670 8240 13740 8260
rect 13670 7080 13680 8240
rect 13720 7080 13740 8240
rect 13670 7060 13740 7080
rect 13770 8240 13850 8260
rect 13770 7080 13790 8240
rect 13830 7080 13850 8240
rect 13770 7060 13850 7080
rect 13880 8240 13960 8260
rect 13880 7080 13900 8240
rect 13940 7080 13960 8240
rect 13880 7060 13960 7080
rect 13990 8240 14070 8260
rect 13990 7080 14010 8240
rect 14050 7080 14070 8240
rect 13990 7060 14070 7080
rect 14100 8240 14180 8260
rect 14100 7080 14120 8240
rect 14160 7080 14180 8240
rect 14100 7060 14180 7080
rect 14210 8240 14290 8260
rect 14210 7080 14230 8240
rect 14270 7080 14290 8240
rect 14210 7060 14290 7080
rect 14320 8240 14400 8260
rect 14320 7080 14340 8240
rect 14380 7080 14400 8240
rect 14320 7060 14400 7080
rect 14430 8240 14510 8260
rect 14430 7080 14450 8240
rect 14490 7080 14510 8240
rect 14430 7060 14510 7080
rect 14540 8240 14620 8260
rect 14540 7080 14560 8240
rect 14600 7080 14620 8240
rect 14540 7060 14620 7080
rect 14650 8240 14730 8260
rect 14650 7080 14670 8240
rect 14710 7080 14730 8240
rect 14650 7060 14730 7080
rect 14760 8240 14840 8260
rect 14760 7080 14780 8240
rect 14820 7080 14840 8240
rect 14760 7060 14840 7080
rect 14870 8240 14950 8260
rect 14870 7080 14890 8240
rect 14930 7080 14950 8240
rect 14870 7060 14950 7080
rect 14980 8240 15060 8260
rect 14980 7080 15000 8240
rect 15040 7080 15060 8240
rect 14980 7060 15060 7080
rect 15090 8240 15170 8260
rect 15090 7080 15110 8240
rect 15150 7080 15170 8240
rect 15090 7060 15170 7080
rect 15200 8240 15280 8260
rect 15200 7080 15220 8240
rect 15260 7080 15280 8240
rect 15200 7060 15280 7080
rect 15310 8240 15390 8260
rect 15310 7080 15330 8240
rect 15370 7080 15390 8240
rect 15310 7060 15390 7080
rect 15420 8240 15500 8260
rect 15420 7080 15440 8240
rect 15480 7080 15500 8240
rect 15420 7060 15500 7080
rect 15530 8240 15610 8260
rect 15530 7080 15550 8240
rect 15590 7080 15610 8240
rect 15530 7060 15610 7080
rect 15640 8240 15720 8260
rect 15640 7080 15660 8240
rect 15700 7080 15720 8240
rect 15640 7060 15720 7080
rect 15750 8240 15830 8260
rect 15750 7080 15770 8240
rect 15810 7080 15830 8240
rect 15750 7060 15830 7080
rect 15860 8240 15940 8260
rect 15860 7080 15880 8240
rect 15920 7080 15940 8240
rect 15860 7060 15940 7080
rect 15970 8240 16050 8260
rect 15970 7080 15990 8240
rect 16030 7080 16050 8240
rect 15970 7060 16050 7080
rect 16080 8240 16160 8260
rect 16080 7080 16100 8240
rect 16140 7080 16160 8240
rect 16080 7060 16160 7080
rect 16190 8240 16270 8260
rect 16190 7080 16210 8240
rect 16250 7080 16270 8240
rect 16190 7060 16270 7080
rect 16300 8240 16380 8260
rect 16300 7080 16320 8240
rect 16360 7080 16380 8240
rect 16300 7060 16380 7080
rect 16410 8240 16490 8260
rect 16410 7080 16430 8240
rect 16470 7080 16490 8240
rect 16410 7060 16490 7080
rect 16520 8240 16600 8260
rect 16520 7080 16540 8240
rect 16580 7080 16600 8240
rect 16520 7060 16600 7080
rect 16630 8240 16710 8260
rect 16630 7080 16650 8240
rect 16690 7080 16710 8240
rect 16630 7060 16710 7080
rect 16740 8240 16820 8260
rect 16740 7080 16760 8240
rect 16800 7080 16820 8240
rect 16740 7060 16820 7080
rect 16850 8240 16930 8260
rect 16850 7080 16870 8240
rect 16910 7080 16930 8240
rect 16850 7060 16930 7080
rect 16960 8240 17030 8260
rect 16960 7080 16980 8240
rect 17020 7080 17030 8240
rect 16960 7060 17030 7080
rect 13630 5840 13700 5860
rect 9870 5600 9940 5620
rect 9870 4440 9880 5600
rect 9920 4440 9940 5600
rect 9870 4420 9940 4440
rect 9970 5600 10050 5620
rect 9970 4440 9990 5600
rect 10030 4440 10050 5600
rect 9970 4420 10050 4440
rect 10080 5600 10160 5620
rect 10080 4440 10100 5600
rect 10140 4440 10160 5600
rect 10080 4420 10160 4440
rect 10190 5600 10270 5620
rect 10190 4440 10210 5600
rect 10250 4440 10270 5600
rect 10190 4420 10270 4440
rect 10300 5600 10380 5620
rect 10300 4440 10320 5600
rect 10360 4440 10380 5600
rect 10300 4420 10380 4440
rect 10410 5600 10490 5620
rect 10410 4440 10430 5600
rect 10470 4440 10490 5600
rect 10410 4420 10490 4440
rect 10520 5600 10600 5620
rect 10520 4440 10540 5600
rect 10580 4440 10600 5600
rect 10520 4420 10600 4440
rect 10630 5600 10710 5620
rect 10630 4440 10650 5600
rect 10690 4440 10710 5600
rect 10630 4420 10710 4440
rect 10740 5600 10820 5620
rect 10740 4440 10760 5600
rect 10800 4440 10820 5600
rect 10740 4420 10820 4440
rect 10850 5600 10930 5620
rect 10850 4440 10870 5600
rect 10910 4440 10930 5600
rect 10850 4420 10930 4440
rect 10960 5600 11040 5620
rect 10960 4440 10980 5600
rect 11020 4440 11040 5600
rect 10960 4420 11040 4440
rect 11070 5600 11150 5620
rect 11070 4440 11090 5600
rect 11130 4440 11150 5600
rect 11070 4420 11150 4440
rect 11180 5600 11260 5620
rect 11180 4440 11200 5600
rect 11240 4440 11260 5600
rect 11180 4420 11260 4440
rect 11290 5600 11370 5620
rect 11290 4440 11310 5600
rect 11350 4440 11370 5600
rect 11290 4420 11370 4440
rect 11400 5600 11480 5620
rect 11400 4440 11420 5600
rect 11460 4440 11480 5600
rect 11400 4420 11480 4440
rect 11510 5600 11590 5620
rect 11510 4440 11530 5600
rect 11570 4440 11590 5600
rect 11510 4420 11590 4440
rect 11620 5600 11700 5620
rect 11620 4440 11640 5600
rect 11680 4440 11700 5600
rect 11620 4420 11700 4440
rect 11730 5600 11810 5620
rect 11730 4440 11750 5600
rect 11790 4440 11810 5600
rect 11730 4420 11810 4440
rect 11840 5600 11920 5620
rect 11840 4440 11860 5600
rect 11900 4440 11920 5600
rect 11840 4420 11920 4440
rect 11950 5600 12030 5620
rect 11950 4440 11970 5600
rect 12010 4440 12030 5600
rect 11950 4420 12030 4440
rect 12060 5600 12140 5620
rect 12060 4440 12080 5600
rect 12120 4440 12140 5600
rect 12060 4420 12140 4440
rect 12170 5600 12250 5620
rect 12170 4440 12190 5600
rect 12230 4440 12250 5600
rect 12170 4420 12250 4440
rect 12280 5600 12360 5620
rect 12280 4440 12300 5600
rect 12340 4440 12360 5600
rect 12280 4420 12360 4440
rect 12390 5600 12470 5620
rect 12390 4440 12410 5600
rect 12450 4440 12470 5600
rect 12390 4420 12470 4440
rect 12500 5600 12580 5620
rect 12500 4440 12520 5600
rect 12560 4440 12580 5600
rect 12500 4420 12580 4440
rect 12610 5600 12690 5620
rect 12610 4440 12630 5600
rect 12670 4440 12690 5600
rect 12610 4420 12690 4440
rect 12720 5600 12800 5620
rect 12720 4440 12740 5600
rect 12780 4440 12800 5600
rect 12720 4420 12800 4440
rect 12830 5600 12910 5620
rect 12830 4440 12850 5600
rect 12890 4440 12910 5600
rect 12830 4420 12910 4440
rect 12940 5600 13020 5620
rect 12940 4440 12960 5600
rect 13000 4440 13020 5600
rect 12940 4420 13020 4440
rect 13050 5600 13130 5620
rect 13050 4440 13070 5600
rect 13110 4440 13130 5600
rect 13050 4420 13130 4440
rect 13160 5600 13230 5620
rect 13160 4440 13180 5600
rect 13220 4440 13230 5600
rect 13630 4680 13640 5840
rect 13680 4680 13700 5840
rect 13630 4660 13700 4680
rect 13730 5840 13810 5860
rect 13730 4680 13750 5840
rect 13790 4680 13810 5840
rect 13730 4660 13810 4680
rect 13840 5840 13920 5860
rect 13840 4680 13860 5840
rect 13900 4680 13920 5840
rect 13840 4660 13920 4680
rect 13950 5840 14030 5860
rect 13950 4680 13970 5840
rect 14010 4680 14030 5840
rect 13950 4660 14030 4680
rect 14060 5840 14140 5860
rect 14060 4680 14080 5840
rect 14120 4680 14140 5840
rect 14060 4660 14140 4680
rect 14170 5840 14250 5860
rect 14170 4680 14190 5840
rect 14230 4680 14250 5840
rect 14170 4660 14250 4680
rect 14280 5840 14360 5860
rect 14280 4680 14300 5840
rect 14340 4680 14360 5840
rect 14280 4660 14360 4680
rect 14390 5840 14470 5860
rect 14390 4680 14410 5840
rect 14450 4680 14470 5840
rect 14390 4660 14470 4680
rect 14500 5840 14580 5860
rect 14500 4680 14520 5840
rect 14560 4680 14580 5840
rect 14500 4660 14580 4680
rect 14610 5840 14690 5860
rect 14610 4680 14630 5840
rect 14670 4680 14690 5840
rect 14610 4660 14690 4680
rect 14720 5840 14800 5860
rect 14720 4680 14740 5840
rect 14780 4680 14800 5840
rect 14720 4660 14800 4680
rect 14830 5840 14910 5860
rect 14830 4680 14850 5840
rect 14890 4680 14910 5840
rect 14830 4660 14910 4680
rect 14940 5840 15020 5860
rect 14940 4680 14960 5840
rect 15000 4680 15020 5840
rect 14940 4660 15020 4680
rect 15050 5840 15130 5860
rect 15050 4680 15070 5840
rect 15110 4680 15130 5840
rect 15050 4660 15130 4680
rect 15160 5840 15240 5860
rect 15160 4680 15180 5840
rect 15220 4680 15240 5840
rect 15160 4660 15240 4680
rect 15270 5840 15350 5860
rect 15270 4680 15290 5840
rect 15330 4680 15350 5840
rect 15270 4660 15350 4680
rect 15380 5840 15460 5860
rect 15380 4680 15400 5840
rect 15440 4680 15460 5840
rect 15380 4660 15460 4680
rect 15490 5840 15570 5860
rect 15490 4680 15510 5840
rect 15550 4680 15570 5840
rect 15490 4660 15570 4680
rect 15600 5840 15680 5860
rect 15600 4680 15620 5840
rect 15660 4680 15680 5840
rect 15600 4660 15680 4680
rect 15710 5840 15790 5860
rect 15710 4680 15730 5840
rect 15770 4680 15790 5840
rect 15710 4660 15790 4680
rect 15820 5840 15900 5860
rect 15820 4680 15840 5840
rect 15880 4680 15900 5840
rect 15820 4660 15900 4680
rect 15930 5840 16010 5860
rect 15930 4680 15950 5840
rect 15990 4680 16010 5840
rect 15930 4660 16010 4680
rect 16040 5840 16120 5860
rect 16040 4680 16060 5840
rect 16100 4680 16120 5840
rect 16040 4660 16120 4680
rect 16150 5840 16230 5860
rect 16150 4680 16170 5840
rect 16210 4680 16230 5840
rect 16150 4660 16230 4680
rect 16260 5840 16340 5860
rect 16260 4680 16280 5840
rect 16320 4680 16340 5840
rect 16260 4660 16340 4680
rect 16370 5840 16450 5860
rect 16370 4680 16390 5840
rect 16430 4680 16450 5840
rect 16370 4660 16450 4680
rect 16480 5840 16560 5860
rect 16480 4680 16500 5840
rect 16540 4680 16560 5840
rect 16480 4660 16560 4680
rect 16590 5840 16670 5860
rect 16590 4680 16610 5840
rect 16650 4680 16670 5840
rect 16590 4660 16670 4680
rect 16700 5840 16780 5860
rect 16700 4680 16720 5840
rect 16760 4680 16780 5840
rect 16700 4660 16780 4680
rect 16810 5840 16890 5860
rect 16810 4680 16830 5840
rect 16870 4680 16890 5840
rect 16810 4660 16890 4680
rect 16920 5840 16990 5860
rect 16920 4680 16940 5840
rect 16980 4680 16990 5840
rect 16920 4660 16990 4680
rect 13160 4420 13230 4440
<< ndiffc >>
rect 23390 41920 23430 42080
rect 21730 41700 21770 41860
rect 21840 41700 21880 41860
rect 23500 41920 23540 42080
rect 22590 41530 22630 41690
rect 22700 41530 22740 41690
rect 22890 41530 22930 41690
rect 23000 41530 23040 41690
rect 23110 41530 23150 41690
rect 23390 41390 23430 41550
rect 23500 41390 23540 41550
rect 5959 41000 5999 41160
rect 6069 41000 6109 41160
rect 6189 41000 6229 41160
rect 6299 41000 6339 41160
rect 6409 41000 6449 41160
rect 6529 41000 6569 41160
rect 6639 41000 6679 41160
rect 6749 41000 6789 41160
rect 6859 41000 6899 41160
rect 6969 41000 7009 41160
rect 7089 41000 7129 41160
rect 7199 41000 7239 41160
rect 7309 41000 7349 41160
rect 7419 41000 7459 41160
rect 7529 41000 7569 41160
rect 7639 41000 7679 41160
rect 7749 41000 7789 41160
rect 7859 41000 7899 41160
rect 7969 41000 8009 41160
rect 8149 41000 8189 41160
rect 8259 41000 8299 41160
rect 8369 41000 8409 41160
rect 8479 41000 8519 41160
rect 8589 41000 8629 41160
rect 8699 41000 8739 41160
rect 8809 41000 8849 41160
rect 8919 41000 8959 41160
rect 9029 41000 9069 41160
rect 9139 41000 9179 41160
rect 9249 41000 9289 41160
rect 9359 41000 9399 41160
rect 9469 41000 9509 41160
rect 9579 41000 9619 41160
rect 9689 41000 9729 41160
rect 9799 41000 9839 41160
rect 9909 41000 9949 41160
rect 2659 39780 2699 40540
rect 2769 39780 2809 40540
rect 2989 39780 3029 40540
rect 3099 39780 3139 40540
rect 6359 39680 6399 39840
rect 6469 39680 6509 39840
rect 6579 39680 6619 39840
rect 6689 39680 6729 39840
rect 6799 39680 6839 39840
rect 6909 39680 6949 39840
rect 7019 39680 7059 39840
rect 7129 39680 7169 39840
rect 7239 39680 7279 39840
rect 7349 39680 7389 39840
rect 7459 39680 7499 39840
rect 7569 39680 7609 39840
rect 7679 39680 7719 39840
rect 7789 39680 7829 39840
rect 7899 39680 7939 39840
rect 8009 39680 8049 39840
rect 8119 39680 8159 39840
rect 8229 39680 8269 39840
rect 8339 39680 8379 39840
rect 8449 39680 8489 39840
rect 8559 39680 8599 39840
rect 8669 39680 8709 39840
rect 8779 39680 8819 39840
rect 8889 39680 8929 39840
rect 8999 39680 9039 39840
rect 9109 39680 9149 39840
rect 9219 39680 9259 39840
rect 9329 39680 9369 39840
rect 9439 39680 9479 39840
rect 9549 39680 9589 39840
rect 9659 39680 9699 39840
rect 9769 39680 9809 39840
rect 9879 39680 9919 39840
rect 3780 36270 3820 37030
rect 3890 36270 3930 37030
rect 4000 36270 4040 37030
rect 4110 36270 4150 37030
rect 4220 36270 4260 37030
rect 4330 36270 4370 37030
rect 4510 36270 4550 37030
rect 4700 36270 4740 37030
rect 4810 36270 4850 37030
rect 4920 36270 4960 37030
rect 5030 36270 5070 37030
rect 5140 36270 5180 37030
rect 5250 36270 5290 37030
rect 5470 36670 5510 37030
rect 5580 36670 5620 37030
rect 5690 36670 5730 37030
rect 5800 36670 5840 37030
rect 5910 36670 5950 37030
rect 6020 36670 6060 37030
rect 6130 36670 6170 37030
rect 6350 36410 6390 36570
rect 6460 36410 6500 36570
rect 6570 36410 6610 36570
rect 6820 36210 6860 36570
rect 7080 36210 7120 36570
rect 7310 36410 7350 36570
rect 7420 36410 7460 36570
rect 7530 36410 7570 36570
rect 7690 36410 7730 36570
rect 7800 36410 7840 36570
rect 7910 36410 7950 36570
rect 8070 36410 8110 36570
rect 8180 36410 8220 36570
rect 8290 36410 8330 36570
rect 8450 36410 8490 36570
rect 8560 36410 8600 36570
rect 8670 36410 8710 36570
rect 8900 36210 8940 36570
rect 9160 36210 9200 36570
rect 9390 36410 9430 36570
rect 9500 36410 9540 36570
rect 9610 36410 9650 36570
rect 9770 36410 9810 36570
rect 9880 36410 9920 36570
rect 9990 36410 10030 36570
rect 10150 36410 10190 36570
rect 10260 36410 10300 36570
rect 10370 36410 10410 36570
rect 10530 36410 10570 36570
rect 10640 36410 10680 36570
rect 10750 36410 10790 36570
rect 16470 35630 16510 35820
rect 16580 35630 16620 35820
rect 16690 35630 16730 35820
rect 16800 35630 16840 35820
rect 16910 35630 16950 35820
rect 17020 35630 17060 35820
rect 17130 35630 17170 35820
rect 16470 34470 16510 35330
rect 16580 34470 16620 35330
rect 16690 34470 16730 35330
rect 16800 34470 16840 35330
rect 16910 34470 16950 35330
rect 17020 34470 17060 35330
rect 17130 34470 17170 35330
rect 17360 34980 17400 35140
rect 17470 34980 17510 35140
rect 17760 34930 17800 35090
rect 17870 34930 17910 35090
rect 18300 34980 18340 35140
rect 18410 34980 18450 35140
rect 18700 34980 18740 35140
rect 18810 34980 18850 35140
rect 19770 34970 19810 35130
rect 19880 34970 19920 35130
rect 20020 34970 20060 35130
rect 20130 34970 20170 35130
rect 21430 35630 21470 35820
rect 21540 35630 21580 35820
rect 21650 35630 21690 35820
rect 21760 35630 21800 35820
rect 21870 35630 21910 35820
rect 21980 35630 22020 35820
rect 22090 35630 22130 35820
rect 17580 34460 17620 34620
rect 17690 34460 17730 34620
rect 18040 34460 18080 34620
rect 18150 34460 18190 34620
rect 18520 34460 18560 34620
rect 18630 34460 18670 34620
rect 18980 34460 19020 34620
rect 19090 34460 19130 34620
rect 19310 34470 19350 34830
rect 19420 34470 19460 34830
rect 19770 34390 19810 34550
rect 19880 34390 19920 34550
rect 21040 34470 21080 34830
rect 21150 34470 21190 34830
rect 21430 34470 21470 35330
rect 21540 34470 21580 35330
rect 21650 34470 21690 35330
rect 21760 34470 21800 35330
rect 21870 34470 21910 35330
rect 21980 34470 22020 35330
rect 22090 34470 22130 35330
rect 22320 34980 22360 35140
rect 22430 34980 22470 35140
rect 22720 34930 22760 35090
rect 22830 34930 22870 35090
rect 23260 34980 23300 35140
rect 23370 34980 23410 35140
rect 23660 34980 23700 35140
rect 23770 34980 23810 35140
rect 24730 34970 24770 35130
rect 24840 34970 24880 35130
rect 24980 34970 25020 35130
rect 25090 34970 25130 35130
rect 22540 34460 22580 34620
rect 22650 34460 22690 34620
rect 23000 34460 23040 34620
rect 23110 34460 23150 34620
rect 23480 34460 23520 34620
rect 23590 34460 23630 34620
rect 23940 34460 23980 34620
rect 24050 34460 24090 34620
rect 24270 34470 24310 34830
rect 24380 34470 24420 34830
rect 24730 34390 24770 34550
rect 24840 34390 24880 34550
rect 2180 30820 2220 31580
rect 2290 30820 2330 31580
rect 2400 30820 2440 31580
rect 2510 30820 2550 31580
rect 2620 30820 2660 31580
rect 2730 30820 2770 31580
rect 2910 30820 2950 31580
rect 3100 30820 3140 31580
rect 3210 30820 3250 31580
rect 3320 30820 3360 31580
rect 3430 30820 3470 31580
rect 3540 30820 3580 31580
rect 3650 30820 3690 31580
rect 3870 31220 3910 31580
rect 3980 31220 4020 31580
rect 4090 31220 4130 31580
rect 4200 31220 4240 31580
rect 4310 31220 4350 31580
rect 4420 31220 4460 31580
rect 4530 31220 4570 31580
rect 4730 31220 4770 31580
rect 4840 31220 4880 31580
rect 4950 31220 4990 31580
rect 5060 31220 5100 31580
rect 5170 31220 5210 31580
rect 5280 31220 5320 31580
rect 5390 31220 5430 31580
rect 5590 31220 5630 31580
rect 5700 31220 5740 31580
rect 5810 31220 5850 31580
rect 5920 31220 5960 31580
rect 6030 31220 6070 31580
rect 6140 31220 6180 31580
rect 6250 31220 6290 31580
rect 14118 31380 14158 31640
rect 14228 31380 14268 31640
rect 16470 31570 16510 31760
rect 16580 31570 16620 31760
rect 16690 31570 16730 31760
rect 16800 31570 16840 31760
rect 16910 31570 16950 31760
rect 17020 31570 17060 31760
rect 17130 31570 17170 31760
rect 6410 31060 6450 31220
rect 6520 31060 6560 31220
rect 6630 31060 6670 31220
rect 6880 30860 6920 31220
rect 7140 30860 7180 31220
rect 7370 31060 7410 31220
rect 7480 31060 7520 31220
rect 7590 31060 7630 31220
rect 7750 31060 7790 31220
rect 7860 31060 7900 31220
rect 7970 31060 8010 31220
rect 8130 31060 8170 31220
rect 8240 31060 8280 31220
rect 8350 31060 8390 31220
rect 8510 31060 8550 31220
rect 8620 31060 8660 31220
rect 8730 31060 8770 31220
rect 8960 30860 9000 31220
rect 9220 30860 9260 31220
rect 9450 31060 9490 31220
rect 9560 31060 9600 31220
rect 9670 31060 9710 31220
rect 9830 31060 9870 31220
rect 9940 31060 9980 31220
rect 10050 31060 10090 31220
rect 10210 31060 10250 31220
rect 10320 31060 10360 31220
rect 10430 31060 10470 31220
rect 10590 31060 10630 31220
rect 10700 31060 10740 31220
rect 10810 31060 10850 31220
rect 10970 31060 11010 31220
rect 11080 31060 11120 31220
rect 11190 31060 11230 31220
rect 16470 30410 16510 31270
rect 16580 30410 16620 31270
rect 16690 30410 16730 31270
rect 16800 30410 16840 31270
rect 16910 30410 16950 31270
rect 17020 30410 17060 31270
rect 17130 30410 17170 31270
rect 17360 30920 17400 31080
rect 17470 30920 17510 31080
rect 17760 30870 17800 31030
rect 17870 30870 17910 31030
rect 18300 30920 18340 31080
rect 18410 30920 18450 31080
rect 18700 30920 18740 31080
rect 18810 30920 18850 31080
rect 20030 30910 20070 31070
rect 20140 30910 20180 31070
rect 20280 30910 20320 31070
rect 20390 30910 20430 31070
rect 21490 31560 21530 31750
rect 21600 31560 21640 31750
rect 21710 31560 21750 31750
rect 21820 31560 21860 31750
rect 21930 31560 21970 31750
rect 22040 31560 22080 31750
rect 22150 31560 22190 31750
rect 17580 30400 17620 30560
rect 17690 30400 17730 30560
rect 18040 30400 18080 30560
rect 18150 30400 18190 30560
rect 18520 30400 18560 30560
rect 18630 30400 18670 30560
rect 18980 30400 19020 30560
rect 19090 30400 19130 30560
rect 19310 30410 19350 30770
rect 19420 30410 19460 30770
rect 19570 30410 19610 30770
rect 19680 30410 19720 30770
rect 20030 30330 20070 30490
rect 20140 30330 20180 30490
rect 21100 30410 21140 30770
rect 21210 30410 21250 30770
rect 21490 30400 21530 31260
rect 21600 30400 21640 31260
rect 21710 30400 21750 31260
rect 21820 30400 21860 31260
rect 21930 30400 21970 31260
rect 22040 30400 22080 31260
rect 22150 30400 22190 31260
rect 22380 30910 22420 31070
rect 22490 30910 22530 31070
rect 22780 30860 22820 31020
rect 22890 30860 22930 31020
rect 23320 30910 23360 31070
rect 23430 30910 23470 31070
rect 23720 30910 23760 31070
rect 23830 30910 23870 31070
rect 24990 30900 25030 31060
rect 25100 30900 25140 31060
rect 25240 30900 25280 31060
rect 25350 30900 25390 31060
rect 22600 30390 22640 30550
rect 22710 30390 22750 30550
rect 23060 30390 23100 30550
rect 23170 30390 23210 30550
rect 23540 30390 23580 30550
rect 23650 30390 23690 30550
rect 24000 30390 24040 30550
rect 24110 30390 24150 30550
rect 24330 30400 24370 30760
rect 24440 30400 24480 30760
rect 24590 30400 24630 30760
rect 24700 30400 24740 30760
rect 24990 30320 25030 30480
rect 25100 30320 25140 30480
rect 7330 24390 7370 24550
rect 7440 24390 7480 24550
rect 7550 24390 7590 24550
rect 7860 24390 7900 24550
rect 7970 24390 8010 24550
rect 8080 24390 8120 24550
rect 8490 24380 8530 24740
rect 8620 24380 8660 24740
rect 8750 24380 8790 24740
rect 8870 24650 8910 24810
rect 8980 24650 9020 24810
rect 9230 24380 9270 24540
rect 9340 24380 9380 24540
rect 9450 24380 9490 24540
rect 9680 24380 9720 24740
rect 9940 24380 9980 24740
rect 10170 24380 10210 24540
rect 10280 24380 10320 24540
rect 10390 24380 10430 24540
rect 10670 24380 10710 24740
rect 10930 24380 10970 24740
rect 11160 24380 11200 24540
rect 11270 24380 11310 24540
rect 11380 24380 11420 24540
rect 11670 24380 11710 24740
rect 11930 24380 11970 24740
rect 12890 24660 12930 24820
rect 13000 24660 13040 24820
rect 13120 24660 13160 24820
rect 13230 24660 13270 24820
rect 13340 24660 13380 24820
rect 13460 24660 13500 24820
rect 13570 24660 13610 24820
rect 13680 24660 13720 24820
rect 13790 24660 13830 24820
rect 13900 24660 13940 24820
rect 14020 24660 14060 24820
rect 14130 24660 14170 24820
rect 14240 24660 14280 24820
rect 14350 24660 14390 24820
rect 14460 24660 14500 24820
rect 14570 24660 14610 24820
rect 14680 24660 14720 24820
rect 14790 24660 14830 24820
rect 14900 24660 14940 24820
rect 15080 24660 15120 24820
rect 15190 24660 15230 24820
rect 15300 24660 15340 24820
rect 15410 24660 15450 24820
rect 15520 24660 15560 24820
rect 15630 24660 15670 24820
rect 15740 24660 15780 24820
rect 15850 24660 15890 24820
rect 15960 24660 16000 24820
rect 16070 24660 16110 24820
rect 16180 24660 16220 24820
rect 16290 24660 16330 24820
rect 16400 24660 16440 24820
rect 16510 24660 16550 24820
rect 16620 24660 16660 24820
rect 16730 24660 16770 24820
rect 16840 24660 16880 24820
rect 17030 24660 17070 24820
rect 17140 24660 17180 24820
rect 17250 24660 17290 24820
rect 17360 24660 17400 24820
rect 17470 24660 17510 24820
rect 17580 24660 17620 24820
rect 17690 24660 17730 24820
rect 17800 24660 17840 24820
rect 17910 24660 17950 24820
rect 18020 24660 18060 24820
rect 18130 24660 18170 24820
rect 18240 24660 18280 24820
rect 18350 24660 18390 24820
rect 18460 24660 18500 24820
rect 18570 24660 18610 24820
rect 18680 24660 18720 24820
rect 18790 24660 18830 24820
rect 18900 24660 18940 24820
rect 19010 24660 19050 24820
rect 19120 24660 19160 24820
rect 19230 24660 19270 24820
rect 19340 24660 19380 24820
rect 19450 24660 19490 24820
rect 19560 24660 19600 24820
rect 19670 24660 19710 24820
rect 19780 24660 19820 24820
rect 19890 24660 19930 24820
rect 20000 24660 20040 24820
rect 20110 24660 20150 24820
rect 20220 24660 20260 24820
rect 20330 24660 20370 24820
rect 20440 24660 20480 24820
rect 20550 24660 20590 24820
rect 12160 24380 12200 24540
rect 12270 24380 12310 24540
rect 12380 24380 12420 24540
rect 12540 24380 12580 24540
rect 12650 24380 12690 24540
rect 12760 24380 12800 24540
rect 7480 22830 7520 23190
rect 7740 22830 7780 23190
rect 7970 23030 8010 23190
rect 8080 23030 8120 23190
rect 8190 23030 8230 23190
rect 8490 22830 8530 23190
rect 8620 22830 8660 23190
rect 8750 22830 8790 23190
rect 9230 23030 9270 23190
rect 9340 23030 9380 23190
rect 9450 23030 9490 23190
rect 8870 22760 8910 22920
rect 8980 22760 9020 22920
rect 9680 22830 9720 23190
rect 9940 22830 9980 23190
rect 10170 23030 10210 23190
rect 10280 23030 10320 23190
rect 10390 23030 10430 23190
rect 10670 22830 10710 23190
rect 10930 22830 10970 23190
rect 11160 23030 11200 23190
rect 11270 23030 11310 23190
rect 11380 23030 11420 23190
rect 11670 22830 11710 23190
rect 11930 22830 11970 23190
rect 12160 23030 12200 23190
rect 12270 23030 12310 23190
rect 12380 23030 12420 23190
rect 12540 23030 12580 23190
rect 12650 23030 12690 23190
rect 12760 23030 12800 23190
rect 12890 22750 12930 22910
rect 13000 22750 13040 22910
rect 13120 22750 13160 22910
rect 13230 22750 13270 22910
rect 13340 22750 13380 22910
rect 13460 22750 13500 22910
rect 13570 22750 13610 22910
rect 13680 22750 13720 22910
rect 13790 22750 13830 22910
rect 13900 22750 13940 22910
rect 14020 22750 14060 22910
rect 14130 22750 14170 22910
rect 14240 22750 14280 22910
rect 14350 22750 14390 22910
rect 14460 22750 14500 22910
rect 14570 22750 14610 22910
rect 14680 22750 14720 22910
rect 14790 22750 14830 22910
rect 14900 22750 14940 22910
rect 15080 22750 15120 22910
rect 15190 22750 15230 22910
rect 15300 22750 15340 22910
rect 15410 22750 15450 22910
rect 15520 22750 15560 22910
rect 15630 22750 15670 22910
rect 15740 22750 15780 22910
rect 15850 22750 15890 22910
rect 15960 22750 16000 22910
rect 16070 22750 16110 22910
rect 16180 22750 16220 22910
rect 16290 22750 16330 22910
rect 16400 22750 16440 22910
rect 16510 22750 16550 22910
rect 16620 22750 16660 22910
rect 16730 22750 16770 22910
rect 16840 22750 16880 22910
rect 17030 22750 17070 22910
rect 17140 22750 17180 22910
rect 17250 22750 17290 22910
rect 17360 22750 17400 22910
rect 17470 22750 17510 22910
rect 17580 22750 17620 22910
rect 17690 22750 17730 22910
rect 17800 22750 17840 22910
rect 17910 22750 17950 22910
rect 18020 22750 18060 22910
rect 18130 22750 18170 22910
rect 18240 22750 18280 22910
rect 18350 22750 18390 22910
rect 18460 22750 18500 22910
rect 18570 22750 18610 22910
rect 18680 22750 18720 22910
rect 18790 22750 18830 22910
rect 18900 22750 18940 22910
rect 19010 22750 19050 22910
rect 19120 22750 19160 22910
rect 19230 22750 19270 22910
rect 19340 22750 19380 22910
rect 19450 22750 19490 22910
rect 19560 22750 19600 22910
rect 19670 22750 19710 22910
rect 19780 22750 19820 22910
rect 19890 22750 19930 22910
rect 20000 22750 20040 22910
rect 20110 22750 20150 22910
rect 20220 22750 20260 22910
rect 20330 22750 20370 22910
rect 20440 22750 20480 22910
rect 20550 22750 20590 22910
rect 7290 17800 7330 17960
rect 7400 17800 7440 17960
rect 7530 17800 7570 17960
rect 7660 17800 7700 17960
rect 7770 17800 7810 17960
rect 7960 17800 8000 17960
rect 8070 17800 8110 17960
rect 8180 17800 8220 17960
rect 8490 17790 8530 18150
rect 8620 17790 8660 18150
rect 8750 17790 8790 18150
rect 8870 18060 8910 18220
rect 8980 18060 9020 18220
rect 9230 17790 9270 17950
rect 9340 17790 9380 17950
rect 9450 17790 9490 17950
rect 9680 17790 9720 18150
rect 9940 17790 9980 18150
rect 10170 17790 10210 17950
rect 10280 17790 10320 17950
rect 10390 17790 10430 17950
rect 10670 17790 10710 18150
rect 10930 17790 10970 18150
rect 11160 17790 11200 17950
rect 11270 17790 11310 17950
rect 11380 17790 11420 17950
rect 11670 17790 11710 18150
rect 11930 17790 11970 18150
rect 12890 18070 12930 18230
rect 13000 18070 13040 18230
rect 13120 18070 13160 18230
rect 13230 18070 13270 18230
rect 13340 18070 13380 18230
rect 13460 18070 13500 18230
rect 13570 18070 13610 18230
rect 13680 18070 13720 18230
rect 13790 18070 13830 18230
rect 13900 18070 13940 18230
rect 14020 18070 14060 18230
rect 14130 18070 14170 18230
rect 14240 18070 14280 18230
rect 14350 18070 14390 18230
rect 14460 18070 14500 18230
rect 14570 18070 14610 18230
rect 14680 18070 14720 18230
rect 14790 18070 14830 18230
rect 14900 18070 14940 18230
rect 15080 18070 15120 18230
rect 15190 18070 15230 18230
rect 15300 18070 15340 18230
rect 15410 18070 15450 18230
rect 15520 18070 15560 18230
rect 15630 18070 15670 18230
rect 15740 18070 15780 18230
rect 15850 18070 15890 18230
rect 15960 18070 16000 18230
rect 16070 18070 16110 18230
rect 16180 18070 16220 18230
rect 16290 18070 16330 18230
rect 16400 18070 16440 18230
rect 16510 18070 16550 18230
rect 16620 18070 16660 18230
rect 16730 18070 16770 18230
rect 16840 18070 16880 18230
rect 17030 18070 17070 18230
rect 17140 18070 17180 18230
rect 17250 18070 17290 18230
rect 17360 18070 17400 18230
rect 17470 18070 17510 18230
rect 17580 18070 17620 18230
rect 17690 18070 17730 18230
rect 17800 18070 17840 18230
rect 17910 18070 17950 18230
rect 18020 18070 18060 18230
rect 18130 18070 18170 18230
rect 18240 18070 18280 18230
rect 18350 18070 18390 18230
rect 18460 18070 18500 18230
rect 18570 18070 18610 18230
rect 18680 18070 18720 18230
rect 18790 18070 18830 18230
rect 18900 18070 18940 18230
rect 19010 18070 19050 18230
rect 19120 18070 19160 18230
rect 19230 18070 19270 18230
rect 19340 18070 19380 18230
rect 19450 18070 19490 18230
rect 19560 18070 19600 18230
rect 19670 18070 19710 18230
rect 19780 18070 19820 18230
rect 19890 18070 19930 18230
rect 20000 18070 20040 18230
rect 20110 18070 20150 18230
rect 20220 18070 20260 18230
rect 20330 18070 20370 18230
rect 20440 18070 20480 18230
rect 20550 18070 20590 18230
rect 12160 17790 12200 17950
rect 12270 17790 12310 17950
rect 12380 17790 12420 17950
rect 12540 17790 12580 17950
rect 12650 17790 12690 17950
rect 12760 17790 12800 17950
rect 9770 15370 9810 15530
rect 9880 15370 9920 15530
rect 9990 15370 10030 15530
rect 10420 15170 10460 15530
rect 10680 15170 10720 15530
rect 10910 15370 10950 15530
rect 11020 15370 11060 15530
rect 11130 15370 11170 15530
rect 11410 15170 11450 15530
rect 11670 15170 11710 15530
rect 11900 15370 11940 15530
rect 12010 15370 12050 15530
rect 12120 15370 12160 15530
rect 12410 15170 12450 15530
rect 12670 15170 12710 15530
rect 12900 15370 12940 15530
rect 13010 15370 13050 15530
rect 13120 15370 13160 15530
rect 13250 15090 13290 15250
rect 13360 15090 13400 15250
rect 13480 15090 13520 15250
rect 13590 15090 13630 15250
rect 13700 15090 13740 15250
rect 13820 15090 13860 15250
rect 13930 15090 13970 15250
rect 14040 15090 14080 15250
rect 14150 15090 14190 15250
rect 14260 15090 14300 15250
rect 14380 15090 14420 15250
rect 14490 15090 14530 15250
rect 14600 15090 14640 15250
rect 14710 15090 14750 15250
rect 14820 15090 14860 15250
rect 14930 15090 14970 15250
rect 15040 15090 15080 15250
rect 15150 15090 15190 15250
rect 15260 15090 15300 15250
rect 15440 15090 15480 15250
rect 15550 15090 15590 15250
rect 15660 15090 15700 15250
rect 15770 15090 15810 15250
rect 15880 15090 15920 15250
rect 15990 15090 16030 15250
rect 16100 15090 16140 15250
rect 16210 15090 16250 15250
rect 16320 15090 16360 15250
rect 16430 15090 16470 15250
rect 16540 15090 16580 15250
rect 16650 15090 16690 15250
rect 16760 15090 16800 15250
rect 16870 15090 16910 15250
rect 16980 15090 17020 15250
rect 17090 15090 17130 15250
rect 17200 15090 17240 15250
rect 17390 15090 17430 15250
rect 17500 15090 17540 15250
rect 17610 15090 17650 15250
rect 17720 15090 17760 15250
rect 17830 15090 17870 15250
rect 17940 15090 17980 15250
rect 18050 15090 18090 15250
rect 18160 15090 18200 15250
rect 18270 15090 18310 15250
rect 18380 15090 18420 15250
rect 18490 15090 18530 15250
rect 18600 15090 18640 15250
rect 18710 15090 18750 15250
rect 18820 15090 18860 15250
rect 18930 15090 18970 15250
rect 19040 15090 19080 15250
rect 19150 15090 19190 15250
rect 19260 15090 19300 15250
rect 19370 15090 19410 15250
rect 19480 15090 19520 15250
rect 19590 15090 19630 15250
rect 19700 15090 19740 15250
rect 19810 15090 19850 15250
rect 19920 15090 19960 15250
rect 20030 15090 20070 15250
rect 20140 15090 20180 15250
rect 20250 15090 20290 15250
rect 20360 15090 20400 15250
rect 20470 15090 20510 15250
rect 20580 15090 20620 15250
rect 20690 15090 20730 15250
rect 20800 15090 20840 15250
rect 20910 15090 20950 15250
rect 7290 12140 7330 12300
rect 7400 12140 7440 12300
rect 7510 12140 7550 12300
rect 7920 12140 7960 12500
rect 8180 12140 8220 12500
rect 8560 12100 8600 12460
rect 8690 12100 8730 12460
rect 8820 12100 8860 12460
rect 8940 12410 8980 12570
rect 9050 12410 9090 12570
rect 9200 12410 9240 12570
rect 9310 12410 9350 12570
rect 9450 12410 9490 12570
rect 9560 12410 9600 12570
rect 9870 12140 9910 12300
rect 9980 12140 10020 12300
rect 10090 12140 10130 12300
rect 10520 12140 10560 12500
rect 10780 12140 10820 12500
rect 11010 12140 11050 12300
rect 11120 12140 11160 12300
rect 11230 12140 11270 12300
rect 11510 12140 11550 12500
rect 11770 12140 11810 12500
rect 12000 12140 12040 12300
rect 12110 12140 12150 12300
rect 12220 12140 12260 12300
rect 12510 12140 12550 12500
rect 12770 12140 12810 12500
rect 13350 12420 13390 12580
rect 13460 12420 13500 12580
rect 13580 12420 13620 12580
rect 13690 12420 13730 12580
rect 13800 12420 13840 12580
rect 13920 12420 13960 12580
rect 14030 12420 14070 12580
rect 14140 12420 14180 12580
rect 14250 12420 14290 12580
rect 14360 12420 14400 12580
rect 14480 12420 14520 12580
rect 14590 12420 14630 12580
rect 14700 12420 14740 12580
rect 14810 12420 14850 12580
rect 14920 12420 14960 12580
rect 15030 12420 15070 12580
rect 15140 12420 15180 12580
rect 15250 12420 15290 12580
rect 15360 12420 15400 12580
rect 15540 12420 15580 12580
rect 15650 12420 15690 12580
rect 15760 12420 15800 12580
rect 15870 12420 15910 12580
rect 15980 12420 16020 12580
rect 16090 12420 16130 12580
rect 16200 12420 16240 12580
rect 16310 12420 16350 12580
rect 16420 12420 16460 12580
rect 16530 12420 16570 12580
rect 16640 12420 16680 12580
rect 16750 12420 16790 12580
rect 16860 12420 16900 12580
rect 16970 12420 17010 12580
rect 17080 12420 17120 12580
rect 17190 12420 17230 12580
rect 17300 12420 17340 12580
rect 17490 12420 17530 12580
rect 17600 12420 17640 12580
rect 17710 12420 17750 12580
rect 17820 12420 17860 12580
rect 17930 12420 17970 12580
rect 18040 12420 18080 12580
rect 18150 12420 18190 12580
rect 18260 12420 18300 12580
rect 18370 12420 18410 12580
rect 18480 12420 18520 12580
rect 18590 12420 18630 12580
rect 18700 12420 18740 12580
rect 18810 12420 18850 12580
rect 18920 12420 18960 12580
rect 19030 12420 19070 12580
rect 19140 12420 19180 12580
rect 19250 12420 19290 12580
rect 19360 12420 19400 12580
rect 19470 12420 19510 12580
rect 19580 12420 19620 12580
rect 19690 12420 19730 12580
rect 19800 12420 19840 12580
rect 19910 12420 19950 12580
rect 20020 12420 20060 12580
rect 20130 12420 20170 12580
rect 20240 12420 20280 12580
rect 20350 12420 20390 12580
rect 20460 12420 20500 12580
rect 20570 12420 20610 12580
rect 20680 12420 20720 12580
rect 20790 12420 20830 12580
rect 20900 12420 20940 12580
rect 21010 12420 21050 12580
rect 13000 12140 13040 12300
rect 13110 12140 13150 12300
rect 13220 12140 13260 12300
rect 7860 11120 7900 11280
rect 7970 11120 8010 11280
rect 8100 11120 8140 11280
rect 8230 11120 8270 11280
rect 8340 11120 8380 11280
rect 7290 10750 7330 10910
rect 7400 10750 7440 10910
rect 7510 10750 7550 10910
rect 8650 10600 8690 10960
rect 8780 10600 8820 10960
rect 8910 10600 8950 10960
rect 9870 10750 9910 10910
rect 9980 10750 10020 10910
rect 10090 10750 10130 10910
rect 9030 10490 9070 10650
rect 9140 10490 9180 10650
rect 9290 10490 9330 10650
rect 9400 10490 9440 10650
rect 9540 10490 9580 10650
rect 9650 10490 9690 10650
rect 10520 10550 10560 10910
rect 10780 10550 10820 10910
rect 11010 10750 11050 10910
rect 11120 10750 11160 10910
rect 11230 10750 11270 10910
rect 11510 10550 11550 10910
rect 11770 10550 11810 10910
rect 12000 10750 12040 10910
rect 12110 10750 12150 10910
rect 12220 10750 12260 10910
rect 12510 10550 12550 10910
rect 12770 10550 12810 10910
rect 13000 10750 13040 10910
rect 13110 10750 13150 10910
rect 13220 10750 13260 10910
rect 13340 10470 13380 10630
rect 13450 10470 13490 10630
rect 13570 10470 13610 10630
rect 13680 10470 13720 10630
rect 13790 10470 13830 10630
rect 13910 10470 13950 10630
rect 14020 10470 14060 10630
rect 14130 10470 14170 10630
rect 14240 10470 14280 10630
rect 14350 10470 14390 10630
rect 14470 10470 14510 10630
rect 14580 10470 14620 10630
rect 14690 10470 14730 10630
rect 14800 10470 14840 10630
rect 14910 10470 14950 10630
rect 15020 10470 15060 10630
rect 15130 10470 15170 10630
rect 15240 10470 15280 10630
rect 15350 10470 15390 10630
rect 15530 10470 15570 10630
rect 15640 10470 15680 10630
rect 15750 10470 15790 10630
rect 15860 10470 15900 10630
rect 15970 10470 16010 10630
rect 16080 10470 16120 10630
rect 16190 10470 16230 10630
rect 16300 10470 16340 10630
rect 16410 10470 16450 10630
rect 16520 10470 16560 10630
rect 16630 10470 16670 10630
rect 16740 10470 16780 10630
rect 16850 10470 16890 10630
rect 16960 10470 17000 10630
rect 17070 10470 17110 10630
rect 17180 10470 17220 10630
rect 17290 10470 17330 10630
rect 17480 10470 17520 10630
rect 17590 10470 17630 10630
rect 17700 10470 17740 10630
rect 17810 10470 17850 10630
rect 17920 10470 17960 10630
rect 18030 10470 18070 10630
rect 18140 10470 18180 10630
rect 18250 10470 18290 10630
rect 18360 10470 18400 10630
rect 18470 10470 18510 10630
rect 18580 10470 18620 10630
rect 18690 10470 18730 10630
rect 18800 10470 18840 10630
rect 18910 10470 18950 10630
rect 19020 10470 19060 10630
rect 19130 10470 19170 10630
rect 19240 10470 19280 10630
rect 19350 10470 19390 10630
rect 19460 10470 19500 10630
rect 19570 10470 19610 10630
rect 19680 10470 19720 10630
rect 19790 10470 19830 10630
rect 19900 10470 19940 10630
rect 20010 10470 20050 10630
rect 20120 10470 20160 10630
rect 20230 10470 20270 10630
rect 20340 10470 20380 10630
rect 20450 10470 20490 10630
rect 20560 10470 20600 10630
rect 20670 10470 20710 10630
rect 20780 10470 20820 10630
rect 20890 10470 20930 10630
rect 21000 10470 21040 10630
rect 9880 3230 9920 3790
rect 9990 3230 10030 3790
rect 10100 3230 10140 3790
rect 10210 3230 10250 3790
rect 10320 3230 10360 3790
rect 10430 3230 10470 3790
rect 10540 3230 10580 3790
rect 10650 3230 10690 3790
rect 10760 3230 10800 3790
rect 10870 3230 10910 3790
rect 10980 3230 11020 3790
rect 11090 3230 11130 3790
rect 11200 3230 11240 3790
rect 11310 3230 11350 3790
rect 11420 3230 11460 3790
rect 11530 3230 11570 3790
rect 11640 3230 11680 3790
rect 11750 3230 11790 3790
rect 11860 3230 11900 3790
rect 11970 3230 12010 3790
rect 12080 3230 12120 3790
rect 12190 3230 12230 3790
rect 12300 3230 12340 3790
rect 12410 3230 12450 3790
rect 12520 3230 12560 3790
rect 12630 3230 12670 3790
rect 12740 3230 12780 3790
rect 12850 3230 12890 3790
rect 12960 3230 13000 3790
rect 13070 3230 13110 3790
rect 13180 3230 13220 3790
rect 13640 3560 13680 4120
rect 13750 3560 13790 4120
rect 13860 3560 13900 4120
rect 13970 3560 14010 4120
rect 14080 3560 14120 4120
rect 14190 3560 14230 4120
rect 14300 3560 14340 4120
rect 14410 3560 14450 4120
rect 14520 3560 14560 4120
rect 14630 3560 14670 4120
rect 14740 3560 14780 4120
rect 14850 3560 14890 4120
rect 14960 3560 15000 4120
rect 15070 3560 15110 4120
rect 15180 3560 15220 4120
rect 15290 3560 15330 4120
rect 15400 3560 15440 4120
rect 15510 3560 15550 4120
rect 15620 3560 15660 4120
rect 15730 3560 15770 4120
rect 15840 3560 15880 4120
rect 15950 3560 15990 4120
rect 16060 3560 16100 4120
rect 16170 3560 16210 4120
rect 16280 3560 16320 4120
rect 16390 3560 16430 4120
rect 16500 3560 16540 4120
rect 16610 3560 16650 4120
rect 16720 3560 16760 4120
rect 16830 3560 16870 4120
rect 16940 3560 16980 4120
rect 24370 2720 25330 2760
rect 24370 2610 25330 2650
rect 24370 2500 25330 2540
rect 24370 2390 25330 2430
rect 24370 2280 25330 2320
rect 24370 2170 25330 2210
rect 24370 2060 25330 2100
rect 9900 750 9940 1310
rect 10010 750 10050 1310
rect 10120 750 10160 1310
rect 10230 750 10270 1310
rect 10340 750 10380 1310
rect 10450 750 10490 1310
rect 10560 750 10600 1310
rect 10670 750 10710 1310
rect 10780 750 10820 1310
rect 10890 750 10930 1310
rect 11000 750 11040 1310
rect 11110 750 11150 1310
rect 11220 750 11260 1310
rect 11330 750 11370 1310
rect 11440 750 11480 1310
rect 11550 750 11590 1310
rect 11660 750 11700 1310
rect 11770 750 11810 1310
rect 11880 750 11920 1310
rect 11990 750 12030 1310
rect 12100 750 12140 1310
rect 12210 750 12250 1310
rect 12320 750 12360 1310
rect 12430 750 12470 1310
rect 12540 750 12580 1310
rect 12650 750 12690 1310
rect 12760 750 12800 1310
rect 12870 750 12910 1310
rect 12980 750 13020 1310
rect 13090 750 13130 1310
rect 13200 750 13240 1310
rect 13640 740 13680 1300
rect 13750 740 13790 1300
rect 13860 740 13900 1300
rect 13970 740 14010 1300
rect 14080 740 14120 1300
rect 14190 740 14230 1300
rect 14300 740 14340 1300
rect 14410 740 14450 1300
rect 14520 740 14560 1300
rect 14630 740 14670 1300
rect 14740 740 14780 1300
rect 14850 740 14890 1300
rect 14960 740 15000 1300
rect 15070 740 15110 1300
rect 15180 740 15220 1300
rect 15290 740 15330 1300
rect 15400 740 15440 1300
rect 15510 740 15550 1300
rect 15620 740 15660 1300
rect 15730 740 15770 1300
rect 15840 740 15880 1300
rect 15950 740 15990 1300
rect 16060 740 16100 1300
rect 16170 740 16210 1300
rect 16280 740 16320 1300
rect 16390 740 16430 1300
rect 16500 740 16540 1300
rect 16610 740 16650 1300
rect 16720 740 16760 1300
rect 16830 740 16870 1300
rect 16940 740 16980 1300
<< pdiffc >>
rect 21730 42200 21770 42860
rect 21840 42200 21880 42860
rect 21960 42200 22000 42860
rect 22070 42200 22110 42860
rect 22590 42210 22630 42870
rect 22700 42210 22740 42870
rect 22890 42210 22930 42870
rect 23000 42210 23040 42870
rect 23110 42210 23150 42870
rect 23470 42500 23510 43160
rect 23580 42500 23620 43160
rect 2569 41740 2609 41900
rect 2679 41740 2719 41900
rect 2789 41740 2829 41900
rect 2899 41740 2939 41900
rect 2449 41020 2489 41380
rect 2559 41020 2599 41380
rect 2669 41020 2709 41380
rect 2779 41020 2819 41380
rect 2889 41020 2929 41380
rect 2999 41020 3039 41380
rect 3399 41090 3439 41800
rect 3509 41090 3549 41800
rect 3619 41090 3659 41800
rect 3729 41090 3769 41800
rect 3839 41090 3879 41800
rect 3949 41090 3989 41800
rect 4059 41090 4099 41800
rect 4169 41090 4209 41800
rect 4279 41090 4319 41800
rect 4549 41080 4589 41790
rect 4659 41080 4699 41790
rect 4769 41080 4809 41790
rect 4879 41080 4919 41790
rect 4989 41080 5029 41790
rect 5099 41080 5139 41790
rect 5209 41080 5249 41790
rect 5319 41080 5359 41790
rect 5429 41080 5469 41790
rect 5959 41360 5999 41820
rect 6069 41360 6109 41820
rect 6189 41360 6229 41820
rect 6299 41360 6339 41820
rect 6409 41360 6449 41820
rect 6529 41360 6569 41820
rect 6639 41360 6679 41820
rect 6749 41360 6789 41820
rect 6859 41360 6899 41820
rect 6969 41360 7009 41820
rect 7089 41360 7129 41820
rect 7199 41360 7239 41820
rect 7309 41360 7349 41820
rect 7419 41360 7459 41820
rect 7529 41360 7569 41820
rect 7639 41360 7679 41820
rect 7749 41360 7789 41820
rect 7859 41360 7899 41820
rect 7969 41360 8009 41820
rect 8149 41360 8189 41820
rect 8259 41360 8299 41820
rect 8369 41360 8409 41820
rect 8479 41360 8519 41820
rect 8589 41360 8629 41820
rect 8699 41360 8739 41820
rect 8809 41360 8849 41820
rect 8919 41360 8959 41820
rect 9029 41360 9069 41820
rect 9139 41360 9179 41820
rect 9249 41360 9289 41820
rect 9359 41360 9399 41820
rect 9469 41360 9509 41820
rect 9579 41360 9619 41820
rect 9689 41360 9729 41820
rect 9799 41360 9839 41820
rect 9909 41360 9949 41820
rect 3269 39800 3309 40510
rect 3379 39800 3419 40510
rect 3489 39800 3529 40510
rect 3599 39800 3639 40510
rect 3709 39800 3749 40510
rect 3819 39800 3859 40510
rect 3929 39800 3969 40510
rect 4039 39800 4079 40510
rect 4149 39800 4189 40510
rect 4549 39800 4589 40510
rect 4659 39800 4699 40510
rect 4769 39800 4809 40510
rect 4879 39800 4919 40510
rect 4989 39800 5029 40510
rect 5099 39800 5139 40510
rect 5209 39800 5249 40510
rect 5319 39800 5359 40510
rect 5429 39800 5469 40510
rect 6359 40040 6399 40500
rect 6469 40040 6509 40500
rect 6579 40040 6619 40500
rect 6689 40040 6729 40500
rect 6799 40040 6839 40500
rect 6909 40040 6949 40500
rect 7019 40040 7059 40500
rect 7129 40040 7169 40500
rect 7239 40040 7279 40500
rect 7349 40040 7389 40500
rect 7459 40040 7499 40500
rect 7569 40040 7609 40500
rect 7679 40040 7719 40500
rect 7789 40040 7829 40500
rect 7899 40040 7939 40500
rect 8009 40040 8049 40500
rect 8119 40040 8159 40500
rect 8229 40040 8269 40500
rect 8339 40040 8379 40500
rect 8449 40040 8489 40500
rect 8559 40040 8599 40500
rect 8669 40040 8709 40500
rect 8779 40040 8819 40500
rect 8889 40040 8929 40500
rect 8999 40040 9039 40500
rect 9109 40040 9149 40500
rect 9219 40040 9259 40500
rect 9329 40040 9369 40500
rect 9439 40040 9479 40500
rect 9549 40040 9589 40500
rect 9659 40040 9699 40500
rect 9769 40040 9809 40500
rect 9879 40040 9919 40500
rect 3780 33710 3820 34670
rect 3890 33710 3930 34670
rect 4000 33710 4040 34670
rect 4110 33710 4150 34670
rect 4220 33710 4260 34670
rect 4330 33710 4370 34670
rect 4510 33710 4560 34670
rect 4700 33710 4740 34670
rect 4810 33710 4850 34670
rect 4920 33710 4960 34670
rect 5030 33710 5070 34670
rect 5140 33710 5180 34670
rect 5250 33710 5290 34670
rect 5470 33780 5510 34740
rect 5580 33780 5620 34740
rect 5690 33780 5730 34740
rect 5800 33780 5840 34740
rect 5910 33780 5950 34740
rect 6020 33780 6060 34740
rect 6130 33780 6170 34740
rect 6350 34280 6390 34740
rect 6460 34280 6500 34740
rect 15350 35790 15390 35950
rect 15460 35790 15500 35950
rect 15570 35790 15610 35950
rect 17470 35600 17510 36060
rect 17580 35600 17620 36060
rect 17720 35600 17760 36060
rect 17830 35600 17870 36060
rect 18040 35600 18080 36060
rect 18150 35600 18190 36060
rect 18410 35600 18450 36060
rect 18520 35600 18560 36060
rect 18660 35600 18700 36060
rect 18770 35600 18810 36060
rect 18980 35600 19020 36060
rect 19090 35600 19130 36060
rect 6570 34280 6610 34740
rect 6820 34270 6860 34730
rect 6950 34270 6990 34730
rect 7080 34270 7120 34730
rect 7310 34270 7350 34730
rect 7420 34270 7460 34730
rect 7530 34270 7570 34730
rect 7690 34270 7730 34730
rect 7800 34270 7840 34730
rect 7910 34270 7950 34730
rect 8070 34270 8110 34730
rect 8180 34270 8220 34730
rect 8290 34270 8330 34730
rect 8450 34270 8490 34730
rect 8560 34270 8600 34730
rect 8670 34270 8710 34730
rect 8900 34270 8940 34730
rect 9030 34270 9070 34730
rect 9160 34270 9200 34730
rect 9390 34270 9430 34730
rect 9500 34270 9540 34730
rect 9610 34270 9650 34730
rect 9770 34270 9810 34730
rect 9880 34270 9920 34730
rect 9990 34270 10030 34730
rect 10150 34270 10190 34730
rect 10260 34270 10300 34730
rect 10370 34270 10410 34730
rect 10530 34270 10570 34730
rect 10640 34270 10680 34730
rect 10750 34270 10790 34730
rect 19310 35030 19350 35990
rect 19420 35030 19460 35990
rect 19770 35620 19810 36080
rect 19880 35620 19920 36080
rect 20020 35620 20060 36080
rect 20130 35620 20170 36080
rect 21040 35030 21080 35990
rect 21150 35030 21190 35990
rect 22430 35600 22470 36060
rect 22540 35600 22580 36060
rect 22680 35600 22720 36060
rect 22790 35600 22830 36060
rect 23000 35600 23040 36060
rect 23110 35600 23150 36060
rect 23370 35600 23410 36060
rect 23480 35600 23520 36060
rect 23620 35600 23660 36060
rect 23730 35600 23770 36060
rect 23940 35600 23980 36060
rect 24050 35600 24090 36060
rect 24270 35030 24310 35990
rect 24380 35030 24420 35990
rect 24730 35620 24770 36080
rect 24840 35620 24880 36080
rect 24980 35620 25020 36080
rect 25090 35620 25130 36080
rect 13898 32060 13938 32220
rect 14008 32060 14048 32220
rect 14118 32060 14158 32220
rect 14228 32060 14268 32220
rect 17470 31540 17510 32000
rect 17580 31540 17620 32000
rect 17720 31540 17760 32000
rect 17830 31540 17870 32000
rect 18040 31540 18080 32000
rect 18150 31540 18190 32000
rect 18410 31540 18450 32000
rect 18520 31540 18560 32000
rect 18660 31540 18700 32000
rect 18770 31540 18810 32000
rect 18980 31540 19020 32000
rect 19090 31540 19130 32000
rect 2180 29460 2220 30420
rect 2290 29460 2330 30420
rect 2400 29460 2440 30420
rect 2510 29460 2550 30420
rect 2620 29460 2660 30420
rect 2730 29460 2770 30420
rect 2910 29460 2960 30420
rect 3100 29460 3140 30420
rect 3210 29460 3250 30420
rect 3320 29460 3360 30420
rect 3430 29460 3470 30420
rect 3540 29460 3580 30420
rect 3650 29460 3690 30420
rect 3870 29530 3910 30490
rect 3980 29530 4020 30490
rect 4090 29530 4130 30490
rect 4200 29530 4240 30490
rect 4310 29530 4350 30490
rect 4420 29530 4460 30490
rect 4530 29530 4570 30490
rect 4730 29530 4770 30490
rect 4840 29530 4880 30490
rect 4950 29530 4990 30490
rect 5060 29530 5100 30490
rect 5170 29530 5210 30490
rect 5280 29530 5320 30490
rect 5390 29530 5430 30490
rect 5590 29530 5630 30490
rect 5700 29530 5740 30490
rect 5810 29530 5850 30490
rect 5920 29530 5960 30490
rect 6030 29530 6070 30490
rect 6140 29530 6180 30490
rect 6250 29530 6290 30490
rect 6410 30130 6450 30590
rect 6520 30130 6560 30590
rect 6630 30130 6670 30590
rect 6880 30120 6920 30580
rect 7010 30120 7050 30580
rect 7140 30120 7180 30580
rect 7370 30120 7410 30580
rect 7480 30120 7520 30580
rect 7590 30120 7630 30580
rect 7750 30120 7790 30580
rect 7860 30120 7900 30580
rect 7970 30120 8010 30580
rect 8130 30120 8170 30580
rect 8240 30120 8280 30580
rect 8350 30120 8390 30580
rect 8510 30120 8550 30580
rect 8620 30120 8660 30580
rect 8730 30120 8770 30580
rect 8960 30120 9000 30580
rect 9090 30120 9130 30580
rect 9220 30120 9260 30580
rect 9450 30120 9490 30580
rect 9560 30120 9600 30580
rect 9670 30120 9710 30580
rect 9830 30120 9870 30580
rect 9940 30120 9980 30580
rect 10050 30120 10090 30580
rect 10210 30120 10250 30580
rect 10320 30120 10360 30580
rect 10430 30120 10470 30580
rect 10590 30120 10630 30580
rect 10700 30120 10740 30580
rect 10810 30120 10850 30580
rect 10970 30120 11010 30580
rect 11080 30120 11120 30580
rect 11190 30120 11230 30580
rect 19310 30970 19350 31930
rect 19420 30970 19460 31930
rect 19570 30970 19610 31930
rect 19680 30970 19720 31930
rect 20030 31540 20070 32000
rect 20140 31540 20180 32000
rect 20280 31540 20320 32000
rect 20390 31540 20430 32000
rect 21100 30970 21140 31930
rect 21210 30970 21250 31930
rect 22490 31530 22530 31990
rect 22600 31530 22640 31990
rect 22740 31530 22780 31990
rect 22850 31530 22890 31990
rect 23060 31530 23100 31990
rect 23170 31530 23210 31990
rect 23430 31530 23470 31990
rect 23540 31530 23580 31990
rect 23680 31530 23720 31990
rect 23790 31530 23830 31990
rect 24000 31530 24040 31990
rect 24110 31530 24150 31990
rect 24330 30960 24370 31920
rect 24440 30960 24480 31920
rect 24590 30960 24630 31920
rect 24700 30960 24740 31920
rect 24990 31550 25030 32010
rect 25100 31550 25140 32010
rect 25240 31550 25280 32010
rect 25350 31550 25390 32010
rect 7330 26010 7370 26470
rect 7440 26010 7480 26470
rect 7550 26010 7590 26470
rect 7860 26010 7900 26470
rect 7970 26010 8010 26470
rect 8080 26010 8120 26470
rect 8490 26020 8530 26480
rect 8620 26020 8660 26480
rect 8750 26020 8790 26480
rect 8870 26020 8910 26480
rect 8980 26020 9020 26480
rect 9230 26020 9270 26480
rect 9340 26020 9380 26480
rect 9450 26020 9490 26480
rect 9680 26020 9720 26480
rect 9810 26020 9850 26480
rect 9940 26020 9980 26480
rect 10170 26020 10210 26480
rect 10280 26020 10320 26480
rect 10390 26020 10430 26480
rect 10670 26020 10710 26480
rect 10800 26020 10840 26480
rect 10930 26020 10970 26480
rect 11160 26020 11200 26480
rect 11270 26020 11310 26480
rect 11380 26020 11420 26480
rect 11670 26020 11710 26480
rect 11800 26020 11840 26480
rect 11930 26020 11970 26480
rect 12160 26020 12200 26480
rect 12270 26020 12310 26480
rect 12380 26020 12420 26480
rect 12540 26020 12580 26480
rect 12650 26020 12690 26480
rect 12760 26020 12800 26480
rect 12890 26020 12930 26480
rect 13000 26020 13040 26480
rect 13120 26020 13160 26480
rect 13230 26020 13270 26480
rect 13340 26020 13380 26480
rect 13460 26020 13500 26480
rect 13570 26020 13610 26480
rect 13680 26020 13720 26480
rect 13790 26020 13830 26480
rect 13900 26020 13940 26480
rect 14020 26020 14060 26480
rect 14130 26020 14170 26480
rect 14240 26020 14280 26480
rect 14350 26020 14390 26480
rect 14460 26020 14500 26480
rect 14570 26020 14610 26480
rect 14680 26020 14720 26480
rect 14790 26020 14830 26480
rect 14900 26020 14940 26480
rect 15080 26020 15120 26480
rect 15190 26020 15230 26480
rect 15300 26020 15340 26480
rect 15410 26020 15450 26480
rect 15520 26020 15560 26480
rect 15630 26020 15670 26480
rect 15740 26020 15780 26480
rect 15850 26020 15890 26480
rect 15960 26020 16000 26480
rect 16070 26020 16110 26480
rect 16180 26020 16220 26480
rect 16290 26020 16330 26480
rect 16400 26020 16440 26480
rect 16510 26020 16550 26480
rect 16620 26020 16660 26480
rect 16730 26020 16770 26480
rect 16840 26020 16880 26480
rect 17030 26020 17070 26480
rect 17140 26020 17180 26480
rect 17250 26020 17290 26480
rect 17360 26020 17400 26480
rect 17470 26020 17510 26480
rect 17580 26020 17620 26480
rect 17690 26020 17730 26480
rect 17800 26020 17840 26480
rect 17910 26020 17950 26480
rect 18020 26020 18060 26480
rect 18130 26020 18170 26480
rect 18240 26020 18280 26480
rect 18350 26020 18390 26480
rect 18460 26020 18500 26480
rect 18570 26020 18610 26480
rect 18680 26020 18720 26480
rect 18790 26020 18830 26480
rect 18900 26020 18940 26480
rect 19010 26020 19050 26480
rect 19120 26020 19160 26480
rect 19230 26020 19270 26480
rect 19340 26020 19380 26480
rect 19450 26020 19490 26480
rect 19560 26020 19600 26480
rect 19670 26020 19710 26480
rect 19780 26020 19820 26480
rect 19890 26020 19930 26480
rect 20000 26020 20040 26480
rect 20110 26020 20150 26480
rect 20220 26020 20260 26480
rect 20330 26020 20370 26480
rect 20440 26020 20480 26480
rect 20550 26020 20590 26480
rect 7480 21100 7520 21560
rect 7610 21100 7650 21560
rect 7740 21100 7780 21560
rect 7970 21100 8010 21560
rect 8080 21100 8120 21560
rect 8190 21100 8230 21560
rect 8490 21090 8530 21550
rect 8620 21090 8660 21550
rect 8750 21090 8790 21550
rect 8870 21090 8910 21550
rect 8980 21090 9020 21550
rect 9230 21090 9270 21550
rect 9340 21090 9380 21550
rect 9450 21090 9490 21550
rect 9680 21090 9720 21550
rect 9810 21090 9850 21550
rect 9940 21090 9980 21550
rect 10170 21090 10210 21550
rect 10280 21090 10320 21550
rect 10390 21090 10430 21550
rect 10670 21090 10710 21550
rect 10800 21090 10840 21550
rect 10930 21090 10970 21550
rect 11160 21090 11200 21550
rect 11270 21090 11310 21550
rect 11380 21090 11420 21550
rect 11670 21090 11710 21550
rect 11800 21090 11840 21550
rect 11930 21090 11970 21550
rect 12160 21090 12200 21550
rect 12270 21090 12310 21550
rect 12380 21090 12420 21550
rect 12540 21090 12580 21550
rect 12650 21090 12690 21550
rect 12760 21090 12800 21550
rect 12890 21090 12930 21550
rect 13000 21090 13040 21550
rect 13120 21090 13160 21550
rect 13230 21090 13270 21550
rect 13340 21090 13380 21550
rect 13460 21090 13500 21550
rect 13570 21090 13610 21550
rect 13680 21090 13720 21550
rect 13790 21090 13830 21550
rect 13900 21090 13940 21550
rect 14020 21090 14060 21550
rect 14130 21090 14170 21550
rect 14240 21090 14280 21550
rect 14350 21090 14390 21550
rect 14460 21090 14500 21550
rect 14570 21090 14610 21550
rect 14680 21090 14720 21550
rect 14790 21090 14830 21550
rect 14900 21090 14940 21550
rect 15080 21090 15120 21550
rect 15190 21090 15230 21550
rect 15300 21090 15340 21550
rect 15410 21090 15450 21550
rect 15520 21090 15560 21550
rect 15630 21090 15670 21550
rect 15740 21090 15780 21550
rect 15850 21090 15890 21550
rect 15960 21090 16000 21550
rect 16070 21090 16110 21550
rect 16180 21090 16220 21550
rect 16290 21090 16330 21550
rect 16400 21090 16440 21550
rect 16510 21090 16550 21550
rect 16620 21090 16660 21550
rect 16730 21090 16770 21550
rect 16840 21090 16880 21550
rect 17030 21090 17070 21550
rect 17140 21090 17180 21550
rect 17250 21090 17290 21550
rect 17360 21090 17400 21550
rect 17470 21090 17510 21550
rect 17580 21090 17620 21550
rect 17690 21090 17730 21550
rect 17800 21090 17840 21550
rect 17910 21090 17950 21550
rect 18020 21090 18060 21550
rect 18130 21090 18170 21550
rect 18240 21090 18280 21550
rect 18350 21090 18390 21550
rect 18460 21090 18500 21550
rect 18570 21090 18610 21550
rect 18680 21090 18720 21550
rect 18790 21090 18830 21550
rect 18900 21090 18940 21550
rect 19010 21090 19050 21550
rect 19120 21090 19160 21550
rect 19230 21090 19270 21550
rect 19340 21090 19380 21550
rect 19450 21090 19490 21550
rect 19560 21090 19600 21550
rect 19670 21090 19710 21550
rect 19780 21090 19820 21550
rect 19890 21090 19930 21550
rect 20000 21090 20040 21550
rect 20110 21090 20150 21550
rect 20220 21090 20260 21550
rect 20330 21090 20370 21550
rect 20440 21090 20480 21550
rect 20550 21090 20590 21550
rect 7400 19380 7440 20340
rect 7660 19380 7700 20340
rect 7960 19880 8000 20340
rect 8070 19880 8110 20340
rect 8180 19880 8220 20340
rect 8490 19430 8530 19890
rect 8620 19430 8660 19890
rect 8750 19430 8790 19890
rect 8870 19430 8910 19890
rect 8980 19430 9020 19890
rect 9230 19430 9270 19890
rect 9340 19430 9380 19890
rect 9450 19430 9490 19890
rect 9680 19430 9720 19890
rect 9810 19430 9850 19890
rect 9940 19430 9980 19890
rect 10170 19430 10210 19890
rect 10280 19430 10320 19890
rect 10390 19430 10430 19890
rect 10670 19430 10710 19890
rect 10800 19430 10840 19890
rect 10930 19430 10970 19890
rect 11160 19430 11200 19890
rect 11270 19430 11310 19890
rect 11380 19430 11420 19890
rect 11670 19430 11710 19890
rect 11800 19430 11840 19890
rect 11930 19430 11970 19890
rect 12160 19430 12200 19890
rect 12270 19430 12310 19890
rect 12380 19430 12420 19890
rect 12540 19430 12580 19890
rect 12650 19430 12690 19890
rect 12760 19430 12800 19890
rect 12890 19430 12930 19890
rect 13000 19430 13040 19890
rect 13120 19430 13160 19890
rect 13230 19430 13270 19890
rect 13340 19430 13380 19890
rect 13460 19430 13500 19890
rect 13570 19430 13610 19890
rect 13680 19430 13720 19890
rect 13790 19430 13830 19890
rect 13900 19430 13940 19890
rect 14020 19430 14060 19890
rect 14130 19430 14170 19890
rect 14240 19430 14280 19890
rect 14350 19430 14390 19890
rect 14460 19430 14500 19890
rect 14570 19430 14610 19890
rect 14680 19430 14720 19890
rect 14790 19430 14830 19890
rect 14900 19430 14940 19890
rect 15080 19430 15120 19890
rect 15190 19430 15230 19890
rect 15300 19430 15340 19890
rect 15410 19430 15450 19890
rect 15520 19430 15560 19890
rect 15630 19430 15670 19890
rect 15740 19430 15780 19890
rect 15850 19430 15890 19890
rect 15960 19430 16000 19890
rect 16070 19430 16110 19890
rect 16180 19430 16220 19890
rect 16290 19430 16330 19890
rect 16400 19430 16440 19890
rect 16510 19430 16550 19890
rect 16620 19430 16660 19890
rect 16730 19430 16770 19890
rect 16840 19430 16880 19890
rect 17030 19430 17070 19890
rect 17140 19430 17180 19890
rect 17250 19430 17290 19890
rect 17360 19430 17400 19890
rect 17470 19430 17510 19890
rect 17580 19430 17620 19890
rect 17690 19430 17730 19890
rect 17800 19430 17840 19890
rect 17910 19430 17950 19890
rect 18020 19430 18060 19890
rect 18130 19430 18170 19890
rect 18240 19430 18280 19890
rect 18350 19430 18390 19890
rect 18460 19430 18500 19890
rect 18570 19430 18610 19890
rect 18680 19430 18720 19890
rect 18790 19430 18830 19890
rect 18900 19430 18940 19890
rect 19010 19430 19050 19890
rect 19120 19430 19160 19890
rect 19230 19430 19270 19890
rect 19340 19430 19380 19890
rect 19450 19430 19490 19890
rect 19560 19430 19600 19890
rect 19670 19430 19710 19890
rect 19780 19430 19820 19890
rect 19890 19430 19930 19890
rect 20000 19430 20040 19890
rect 20110 19430 20150 19890
rect 20220 19430 20260 19890
rect 20330 19430 20370 19890
rect 20440 19430 20480 19890
rect 20550 19430 20590 19890
rect 9770 14430 9810 14890
rect 9880 14430 9920 14890
rect 9990 14430 10030 14890
rect 10420 14430 10460 14890
rect 10550 14430 10590 14890
rect 10680 14430 10720 14890
rect 10910 14430 10950 14890
rect 11020 14430 11060 14890
rect 11130 14430 11170 14890
rect 11410 14430 11450 14890
rect 11540 14430 11580 14890
rect 11670 14430 11710 14890
rect 11900 14430 11940 14890
rect 12010 14430 12050 14890
rect 12120 14430 12160 14890
rect 12410 14430 12450 14890
rect 12540 14430 12580 14890
rect 12670 14430 12710 14890
rect 12900 14430 12940 14890
rect 13010 14430 13050 14890
rect 13120 14430 13160 14890
rect 13250 14430 13290 14890
rect 13360 14430 13400 14890
rect 13480 14430 13520 14890
rect 13590 14430 13630 14890
rect 13700 14430 13740 14890
rect 13820 14430 13860 14890
rect 13930 14430 13970 14890
rect 14040 14430 14080 14890
rect 14150 14430 14190 14890
rect 14260 14430 14300 14890
rect 14380 14430 14420 14890
rect 14490 14430 14530 14890
rect 14600 14430 14640 14890
rect 14710 14430 14750 14890
rect 14820 14430 14860 14890
rect 14930 14430 14970 14890
rect 15040 14430 15080 14890
rect 15150 14430 15190 14890
rect 15260 14430 15300 14890
rect 15440 14430 15480 14890
rect 15550 14430 15590 14890
rect 15660 14430 15700 14890
rect 15770 14430 15810 14890
rect 15880 14430 15920 14890
rect 15990 14430 16030 14890
rect 16100 14430 16140 14890
rect 16210 14430 16250 14890
rect 16320 14430 16360 14890
rect 16430 14430 16470 14890
rect 16540 14430 16580 14890
rect 16650 14430 16690 14890
rect 16760 14430 16800 14890
rect 16870 14430 16910 14890
rect 16980 14430 17020 14890
rect 17090 14430 17130 14890
rect 17200 14430 17240 14890
rect 17390 14430 17430 14890
rect 17500 14430 17540 14890
rect 17610 14430 17650 14890
rect 17720 14430 17760 14890
rect 17830 14430 17870 14890
rect 17940 14430 17980 14890
rect 18050 14430 18090 14890
rect 18160 14430 18200 14890
rect 18270 14430 18310 14890
rect 18380 14430 18420 14890
rect 18490 14430 18530 14890
rect 18600 14430 18640 14890
rect 18710 14430 18750 14890
rect 18820 14430 18860 14890
rect 18930 14430 18970 14890
rect 19040 14430 19080 14890
rect 19150 14430 19190 14890
rect 19260 14430 19300 14890
rect 19370 14430 19410 14890
rect 19480 14430 19520 14890
rect 19590 14430 19630 14890
rect 19700 14430 19740 14890
rect 19810 14430 19850 14890
rect 19920 14430 19960 14890
rect 20030 14430 20070 14890
rect 20140 14430 20180 14890
rect 20250 14430 20290 14890
rect 20360 14430 20400 14890
rect 20470 14430 20510 14890
rect 20580 14430 20620 14890
rect 20690 14430 20730 14890
rect 20800 14430 20840 14890
rect 20910 14430 20950 14890
rect 7290 12780 7330 13240
rect 7400 12780 7440 13240
rect 7510 12780 7550 13240
rect 7920 12780 7960 13240
rect 8050 12780 8090 13240
rect 8180 12780 8220 13240
rect 8560 12780 8600 13240
rect 8690 12780 8730 13240
rect 8820 12780 8860 13240
rect 8940 12780 8980 13240
rect 9050 12780 9090 13240
rect 9200 12780 9240 13240
rect 9310 12780 9350 13240
rect 9450 12780 9490 13240
rect 9560 12780 9600 13240
rect 9870 12780 9910 13240
rect 9980 12780 10020 13240
rect 10090 12780 10130 13240
rect 10520 12780 10560 13240
rect 10650 12780 10690 13240
rect 10780 12780 10820 13240
rect 11010 12780 11050 13240
rect 11120 12780 11160 13240
rect 11230 12780 11270 13240
rect 11510 12780 11550 13240
rect 11640 12780 11680 13240
rect 11770 12780 11810 13240
rect 12000 12780 12040 13240
rect 12110 12780 12150 13240
rect 12220 12780 12260 13240
rect 12510 12780 12550 13240
rect 12640 12780 12680 13240
rect 12770 12780 12810 13240
rect 13000 12780 13040 13240
rect 13110 12780 13150 13240
rect 13220 12780 13260 13240
rect 13350 12780 13390 13240
rect 13460 12780 13500 13240
rect 13580 12780 13620 13240
rect 13690 12780 13730 13240
rect 13800 12780 13840 13240
rect 13920 12780 13960 13240
rect 14030 12780 14070 13240
rect 14140 12780 14180 13240
rect 14250 12780 14290 13240
rect 14360 12780 14400 13240
rect 14480 12780 14520 13240
rect 14590 12780 14630 13240
rect 14700 12780 14740 13240
rect 14810 12780 14850 13240
rect 14920 12780 14960 13240
rect 15030 12780 15070 13240
rect 15140 12780 15180 13240
rect 15250 12780 15290 13240
rect 15360 12780 15400 13240
rect 15540 12780 15580 13240
rect 15650 12780 15690 13240
rect 15760 12780 15800 13240
rect 15870 12780 15910 13240
rect 15980 12780 16020 13240
rect 16090 12780 16130 13240
rect 16200 12780 16240 13240
rect 16310 12780 16350 13240
rect 16420 12780 16460 13240
rect 16530 12780 16570 13240
rect 16640 12780 16680 13240
rect 16750 12780 16790 13240
rect 16860 12780 16900 13240
rect 16970 12780 17010 13240
rect 17080 12780 17120 13240
rect 17190 12780 17230 13240
rect 17300 12780 17340 13240
rect 17490 12780 17530 13240
rect 17600 12780 17640 13240
rect 17710 12780 17750 13240
rect 17820 12780 17860 13240
rect 17930 12780 17970 13240
rect 18040 12780 18080 13240
rect 18150 12780 18190 13240
rect 18260 12780 18300 13240
rect 18370 12780 18410 13240
rect 18480 12780 18520 13240
rect 18590 12780 18630 13240
rect 18700 12780 18740 13240
rect 18810 12780 18850 13240
rect 18920 12780 18960 13240
rect 19030 12780 19070 13240
rect 19140 12780 19180 13240
rect 19250 12780 19290 13240
rect 19360 12780 19400 13240
rect 19470 12780 19510 13240
rect 19580 12780 19620 13240
rect 19690 12780 19730 13240
rect 19800 12780 19840 13240
rect 19910 12780 19950 13240
rect 20020 12780 20060 13240
rect 20130 12780 20170 13240
rect 20240 12780 20280 13240
rect 20350 12780 20390 13240
rect 20460 12780 20500 13240
rect 20570 12780 20610 13240
rect 20680 12780 20720 13240
rect 20790 12780 20830 13240
rect 20900 12780 20940 13240
rect 21010 12780 21050 13240
rect 7290 9810 7330 10270
rect 7400 9810 7440 10270
rect 7510 9810 7550 10270
rect 7970 9740 8010 10700
rect 8230 9740 8270 10700
rect 8650 9820 8690 10280
rect 8780 9820 8820 10280
rect 8910 9820 8950 10280
rect 9030 9820 9070 10280
rect 9140 9820 9180 10280
rect 9290 9820 9330 10280
rect 9400 9820 9440 10280
rect 9540 9820 9580 10280
rect 9650 9820 9690 10280
rect 9870 9810 9910 10270
rect 9980 9810 10020 10270
rect 10090 9810 10130 10270
rect 10520 9810 10560 10270
rect 10650 9810 10690 10270
rect 10780 9810 10820 10270
rect 11010 9810 11050 10270
rect 11120 9810 11160 10270
rect 11230 9810 11270 10270
rect 11510 9810 11550 10270
rect 11640 9810 11680 10270
rect 11770 9810 11810 10270
rect 12000 9810 12040 10270
rect 12110 9810 12150 10270
rect 12220 9810 12260 10270
rect 12510 9810 12550 10270
rect 12640 9810 12680 10270
rect 12770 9810 12810 10270
rect 13000 9810 13040 10270
rect 13110 9810 13150 10270
rect 13220 9810 13260 10270
rect 13340 9810 13380 10270
rect 13450 9810 13490 10270
rect 13570 9810 13610 10270
rect 13680 9810 13720 10270
rect 13790 9810 13830 10270
rect 13910 9810 13950 10270
rect 14020 9810 14060 10270
rect 14130 9810 14170 10270
rect 14240 9810 14280 10270
rect 14350 9810 14390 10270
rect 14470 9810 14510 10270
rect 14580 9810 14620 10270
rect 14690 9810 14730 10270
rect 14800 9810 14840 10270
rect 14910 9810 14950 10270
rect 15020 9810 15060 10270
rect 15130 9810 15170 10270
rect 15240 9810 15280 10270
rect 15350 9810 15390 10270
rect 15530 9810 15570 10270
rect 15640 9810 15680 10270
rect 15750 9810 15790 10270
rect 15860 9810 15900 10270
rect 15970 9810 16010 10270
rect 16080 9810 16120 10270
rect 16190 9810 16230 10270
rect 16300 9810 16340 10270
rect 16410 9810 16450 10270
rect 16520 9810 16560 10270
rect 16630 9810 16670 10270
rect 16740 9810 16780 10270
rect 16850 9810 16890 10270
rect 16960 9810 17000 10270
rect 17070 9810 17110 10270
rect 17180 9810 17220 10270
rect 17290 9810 17330 10270
rect 17480 9810 17520 10270
rect 17590 9810 17630 10270
rect 17700 9810 17740 10270
rect 17810 9810 17850 10270
rect 17920 9810 17960 10270
rect 18030 9810 18070 10270
rect 18140 9810 18180 10270
rect 18250 9810 18290 10270
rect 18360 9810 18400 10270
rect 18470 9810 18510 10270
rect 18580 9810 18620 10270
rect 18690 9810 18730 10270
rect 18800 9810 18840 10270
rect 18910 9810 18950 10270
rect 19020 9810 19060 10270
rect 19130 9810 19170 10270
rect 19240 9810 19280 10270
rect 19350 9810 19390 10270
rect 19460 9810 19500 10270
rect 19570 9810 19610 10270
rect 19680 9810 19720 10270
rect 19790 9810 19830 10270
rect 19900 9810 19940 10270
rect 20010 9810 20050 10270
rect 20120 9810 20160 10270
rect 20230 9810 20270 10270
rect 20340 9810 20380 10270
rect 20450 9810 20490 10270
rect 20560 9810 20600 10270
rect 20670 9810 20710 10270
rect 20780 9810 20820 10270
rect 20890 9810 20930 10270
rect 21000 9810 21040 10270
rect 9910 7080 9950 8240
rect 10020 7080 10060 8240
rect 10130 7080 10170 8240
rect 10240 7080 10280 8240
rect 10350 7080 10390 8240
rect 10460 7080 10500 8240
rect 10570 7080 10610 8240
rect 10680 7080 10720 8240
rect 10790 7080 10830 8240
rect 10900 7080 10940 8240
rect 11010 7080 11050 8240
rect 11120 7080 11160 8240
rect 11230 7080 11270 8240
rect 11340 7080 11380 8240
rect 11450 7080 11490 8240
rect 11560 7080 11600 8240
rect 11670 7080 11710 8240
rect 11780 7080 11820 8240
rect 11890 7080 11930 8240
rect 12000 7080 12040 8240
rect 12110 7080 12150 8240
rect 12220 7080 12260 8240
rect 12330 7080 12370 8240
rect 12440 7080 12480 8240
rect 12550 7080 12590 8240
rect 12660 7080 12700 8240
rect 12770 7080 12810 8240
rect 12880 7080 12920 8240
rect 12990 7080 13030 8240
rect 13100 7080 13140 8240
rect 13210 7080 13250 8240
rect 13680 7080 13720 8240
rect 13790 7080 13830 8240
rect 13900 7080 13940 8240
rect 14010 7080 14050 8240
rect 14120 7080 14160 8240
rect 14230 7080 14270 8240
rect 14340 7080 14380 8240
rect 14450 7080 14490 8240
rect 14560 7080 14600 8240
rect 14670 7080 14710 8240
rect 14780 7080 14820 8240
rect 14890 7080 14930 8240
rect 15000 7080 15040 8240
rect 15110 7080 15150 8240
rect 15220 7080 15260 8240
rect 15330 7080 15370 8240
rect 15440 7080 15480 8240
rect 15550 7080 15590 8240
rect 15660 7080 15700 8240
rect 15770 7080 15810 8240
rect 15880 7080 15920 8240
rect 15990 7080 16030 8240
rect 16100 7080 16140 8240
rect 16210 7080 16250 8240
rect 16320 7080 16360 8240
rect 16430 7080 16470 8240
rect 16540 7080 16580 8240
rect 16650 7080 16690 8240
rect 16760 7080 16800 8240
rect 16870 7080 16910 8240
rect 16980 7080 17020 8240
rect 9880 4440 9920 5600
rect 9990 4440 10030 5600
rect 10100 4440 10140 5600
rect 10210 4440 10250 5600
rect 10320 4440 10360 5600
rect 10430 4440 10470 5600
rect 10540 4440 10580 5600
rect 10650 4440 10690 5600
rect 10760 4440 10800 5600
rect 10870 4440 10910 5600
rect 10980 4440 11020 5600
rect 11090 4440 11130 5600
rect 11200 4440 11240 5600
rect 11310 4440 11350 5600
rect 11420 4440 11460 5600
rect 11530 4440 11570 5600
rect 11640 4440 11680 5600
rect 11750 4440 11790 5600
rect 11860 4440 11900 5600
rect 11970 4440 12010 5600
rect 12080 4440 12120 5600
rect 12190 4440 12230 5600
rect 12300 4440 12340 5600
rect 12410 4440 12450 5600
rect 12520 4440 12560 5600
rect 12630 4440 12670 5600
rect 12740 4440 12780 5600
rect 12850 4440 12890 5600
rect 12960 4440 13000 5600
rect 13070 4440 13110 5600
rect 13180 4440 13220 5600
rect 13640 4680 13680 5840
rect 13750 4680 13790 5840
rect 13860 4680 13900 5840
rect 13970 4680 14010 5840
rect 14080 4680 14120 5840
rect 14190 4680 14230 5840
rect 14300 4680 14340 5840
rect 14410 4680 14450 5840
rect 14520 4680 14560 5840
rect 14630 4680 14670 5840
rect 14740 4680 14780 5840
rect 14850 4680 14890 5840
rect 14960 4680 15000 5840
rect 15070 4680 15110 5840
rect 15180 4680 15220 5840
rect 15290 4680 15330 5840
rect 15400 4680 15440 5840
rect 15510 4680 15550 5840
rect 15620 4680 15660 5840
rect 15730 4680 15770 5840
rect 15840 4680 15880 5840
rect 15950 4680 15990 5840
rect 16060 4680 16100 5840
rect 16170 4680 16210 5840
rect 16280 4680 16320 5840
rect 16390 4680 16430 5840
rect 16500 4680 16540 5840
rect 16610 4680 16650 5840
rect 16720 4680 16760 5840
rect 16830 4680 16870 5840
rect 16940 4680 16980 5840
<< psubdiff >>
rect 3049 41680 3209 41700
rect 3049 41640 3089 41680
rect 3169 41640 3209 41680
rect 3049 41620 3209 41640
rect 21590 41160 23630 41180
rect 21590 41090 21620 41160
rect 21680 41090 21720 41160
rect 21780 41090 21830 41160
rect 21890 41090 21930 41160
rect 21990 41090 22030 41160
rect 22090 41090 22130 41160
rect 22190 41090 22230 41160
rect 22290 41090 22330 41160
rect 22390 41090 22430 41160
rect 22490 41090 22530 41160
rect 22590 41090 22630 41160
rect 22690 41090 22730 41160
rect 22790 41090 22830 41160
rect 22890 41090 22930 41160
rect 22990 41090 23030 41160
rect 23090 41090 23130 41160
rect 23190 41090 23230 41160
rect 23290 41090 23330 41160
rect 23390 41090 23430 41160
rect 23490 41090 23530 41160
rect 23590 41090 23630 41160
rect 21590 41080 23630 41090
rect 5949 40910 9979 40920
rect 5949 40850 6009 40910
rect 6070 40850 9979 40910
rect 5949 40840 9979 40850
rect 2619 39560 9979 39570
rect 2619 39500 2649 39560
rect 2709 39500 2749 39560
rect 2809 39500 2849 39560
rect 2909 39500 2949 39560
rect 3009 39500 3049 39560
rect 3109 39500 3149 39560
rect 3209 39500 3249 39560
rect 3309 39500 3349 39560
rect 3409 39500 3449 39560
rect 3509 39500 3549 39560
rect 3609 39500 3649 39560
rect 3709 39500 3749 39560
rect 3809 39500 3849 39560
rect 3909 39500 3949 39560
rect 4009 39500 4049 39560
rect 4109 39500 4149 39560
rect 4209 39500 4249 39560
rect 4309 39500 4349 39560
rect 4409 39500 4449 39560
rect 4509 39500 4549 39560
rect 4609 39500 4649 39560
rect 4709 39500 4749 39560
rect 4809 39500 4849 39560
rect 4909 39500 4949 39560
rect 5009 39500 5049 39560
rect 5109 39500 5149 39560
rect 5209 39500 5249 39560
rect 5309 39500 6349 39560
rect 6409 39500 6449 39560
rect 6509 39500 6549 39560
rect 6609 39500 6649 39560
rect 6709 39500 6749 39560
rect 6809 39500 6849 39560
rect 6909 39500 6949 39560
rect 7009 39500 7049 39560
rect 7109 39500 7149 39560
rect 7209 39500 7249 39560
rect 7309 39500 7349 39560
rect 7409 39500 7479 39560
rect 7539 39500 7579 39560
rect 7639 39500 7679 39560
rect 7739 39500 7779 39560
rect 7839 39500 7879 39560
rect 7939 39500 7979 39560
rect 8039 39500 8079 39560
rect 8139 39500 8179 39560
rect 8239 39500 8279 39560
rect 8339 39500 8379 39560
rect 8439 39500 8479 39560
rect 8539 39500 8629 39560
rect 8689 39500 8729 39560
rect 8789 39500 8829 39560
rect 8889 39500 8929 39560
rect 8989 39500 9029 39560
rect 9089 39500 9129 39560
rect 9189 39500 9229 39560
rect 9289 39500 9329 39560
rect 9389 39500 9429 39560
rect 9489 39500 9529 39560
rect 9589 39500 9629 39560
rect 9689 39500 9739 39560
rect 9799 39500 9839 39560
rect 9899 39500 9979 39560
rect 2619 39490 9979 39500
rect 3770 37180 6200 37190
rect 3770 37120 3810 37180
rect 3870 37120 3910 37180
rect 3970 37120 4010 37180
rect 4070 37120 4110 37180
rect 4170 37120 4210 37180
rect 4270 37120 4310 37180
rect 4370 37120 4410 37180
rect 4470 37120 4510 37180
rect 4570 37120 4610 37180
rect 4670 37120 4710 37180
rect 4770 37120 4810 37180
rect 4870 37120 4910 37180
rect 4970 37120 5010 37180
rect 5070 37120 5110 37180
rect 5170 37120 5210 37180
rect 5270 37120 5310 37180
rect 5370 37120 5410 37180
rect 5470 37120 5510 37180
rect 5570 37120 5610 37180
rect 5670 37120 5710 37180
rect 5770 37120 5810 37180
rect 5870 37120 5910 37180
rect 5970 37120 6010 37180
rect 6070 37120 6110 37180
rect 6170 37120 6200 37180
rect 3770 37110 6200 37120
rect 6340 36720 10880 36730
rect 6340 36660 6380 36720
rect 6440 36660 6480 36720
rect 6540 36660 6580 36720
rect 6640 36660 6680 36720
rect 6740 36660 6780 36720
rect 6840 36660 6880 36720
rect 6940 36660 6980 36720
rect 7040 36660 7080 36720
rect 7140 36660 7180 36720
rect 7240 36660 7280 36720
rect 7340 36660 7380 36720
rect 7440 36660 7480 36720
rect 7540 36660 7580 36720
rect 7640 36660 7680 36720
rect 7740 36660 7780 36720
rect 7840 36660 7880 36720
rect 7940 36660 7980 36720
rect 8040 36660 8080 36720
rect 8140 36660 8180 36720
rect 8240 36660 8280 36720
rect 8340 36660 8380 36720
rect 8440 36660 8480 36720
rect 8540 36660 8580 36720
rect 8640 36660 8680 36720
rect 8740 36660 8780 36720
rect 8840 36660 8880 36720
rect 8940 36660 8980 36720
rect 9040 36660 9080 36720
rect 9140 36660 9180 36720
rect 9240 36660 9280 36720
rect 9340 36660 9380 36720
rect 9440 36660 9480 36720
rect 9540 36660 9580 36720
rect 9640 36660 9680 36720
rect 9740 36660 9780 36720
rect 9840 36660 9880 36720
rect 9940 36660 9980 36720
rect 10040 36660 10080 36720
rect 10140 36660 10180 36720
rect 10240 36660 10280 36720
rect 10340 36660 10380 36720
rect 10440 36660 10480 36720
rect 10540 36660 10580 36720
rect 10640 36660 10680 36720
rect 10740 36660 10780 36720
rect 10840 36660 10880 36720
rect 6340 36650 10880 36660
rect 15760 35630 15930 35640
rect 15760 35570 15790 35630
rect 15900 35570 15930 35630
rect 15760 35560 15930 35570
rect 16460 34200 25450 34210
rect 16460 34130 16510 34200
rect 16570 34130 16610 34200
rect 16670 34130 16710 34200
rect 16770 34130 16810 34200
rect 16870 34130 16910 34200
rect 16970 34130 17010 34200
rect 17070 34130 17110 34200
rect 17170 34130 17210 34200
rect 17270 34130 17310 34200
rect 17370 34130 17410 34200
rect 17470 34130 17510 34200
rect 17570 34130 17610 34200
rect 17670 34130 17710 34200
rect 17770 34130 17810 34200
rect 17870 34130 17910 34200
rect 17970 34130 18010 34200
rect 18070 34130 18110 34200
rect 18170 34130 18210 34200
rect 18270 34130 18310 34200
rect 18370 34130 18410 34200
rect 18470 34130 18510 34200
rect 18570 34130 18610 34200
rect 18670 34130 18710 34200
rect 18770 34130 18810 34200
rect 18870 34130 18910 34200
rect 18970 34130 19010 34200
rect 19070 34130 19110 34200
rect 19170 34130 19210 34200
rect 19270 34130 19310 34200
rect 19370 34130 19410 34200
rect 19470 34130 19510 34200
rect 19570 34130 19610 34200
rect 19670 34130 19710 34200
rect 19770 34130 19810 34200
rect 19870 34130 19910 34200
rect 19970 34130 20010 34200
rect 20070 34130 20110 34200
rect 20170 34130 20210 34200
rect 20270 34130 20310 34200
rect 20370 34130 20410 34200
rect 20470 34130 20510 34200
rect 20570 34130 20610 34200
rect 20670 34130 20710 34200
rect 20770 34130 20810 34200
rect 20870 34130 20910 34200
rect 20970 34130 21010 34200
rect 21070 34130 21110 34200
rect 21170 34130 21210 34200
rect 21270 34130 21310 34200
rect 21370 34130 21410 34200
rect 21470 34130 21510 34200
rect 21570 34130 21610 34200
rect 21670 34130 21710 34200
rect 21770 34130 21810 34200
rect 21870 34130 21910 34200
rect 21970 34130 22010 34200
rect 22070 34130 22110 34200
rect 22170 34130 22210 34200
rect 22270 34130 22310 34200
rect 22370 34130 22410 34200
rect 22470 34130 22510 34200
rect 22570 34130 22610 34200
rect 22670 34130 22710 34200
rect 22770 34130 22810 34200
rect 22870 34130 22910 34200
rect 22970 34130 23010 34200
rect 23070 34130 23110 34200
rect 23170 34130 23210 34200
rect 23270 34130 23310 34200
rect 23370 34130 23410 34200
rect 23470 34130 23510 34200
rect 23570 34130 23620 34200
rect 23680 34130 23720 34200
rect 23780 34130 23820 34200
rect 23880 34130 23920 34200
rect 23980 34130 24020 34200
rect 24080 34130 24120 34200
rect 24180 34130 24220 34200
rect 24280 34130 24320 34200
rect 24380 34130 24420 34200
rect 24480 34130 24520 34200
rect 24580 34130 24620 34200
rect 24680 34130 24720 34200
rect 24780 34130 24820 34200
rect 24880 34130 24920 34200
rect 24980 34130 25020 34200
rect 25080 34130 25120 34200
rect 25180 34130 25220 34200
rect 25280 34130 25320 34200
rect 25380 34130 25450 34200
rect 16460 34120 25450 34130
rect 14370 32010 14540 32020
rect 14370 31950 14400 32010
rect 14510 31950 14540 32010
rect 14370 31940 14540 31950
rect 2170 31730 6310 31740
rect 2170 31670 2210 31730
rect 2270 31670 2310 31730
rect 2370 31670 2410 31730
rect 2470 31670 2510 31730
rect 2570 31670 2610 31730
rect 2670 31670 2710 31730
rect 2770 31670 2810 31730
rect 2870 31670 2910 31730
rect 2970 31670 3010 31730
rect 3070 31670 3110 31730
rect 3170 31670 3210 31730
rect 3270 31670 3310 31730
rect 3370 31670 3410 31730
rect 3470 31670 3510 31730
rect 3570 31670 3610 31730
rect 3670 31670 3710 31730
rect 3770 31670 3810 31730
rect 3870 31670 3910 31730
rect 3970 31670 4010 31730
rect 4070 31670 4110 31730
rect 4170 31670 4210 31730
rect 4270 31670 4310 31730
rect 4370 31670 4410 31730
rect 4470 31670 4510 31730
rect 4570 31670 4610 31730
rect 4670 31670 4710 31730
rect 4770 31670 4810 31730
rect 4870 31670 4910 31730
rect 4970 31670 5010 31730
rect 5070 31670 5110 31730
rect 5170 31670 5210 31730
rect 5270 31670 5310 31730
rect 5370 31670 5410 31730
rect 5470 31670 5510 31730
rect 5570 31670 5610 31730
rect 5670 31670 5710 31730
rect 5770 31670 5810 31730
rect 5870 31670 5910 31730
rect 5970 31670 6010 31730
rect 6070 31670 6110 31730
rect 6170 31670 6210 31730
rect 6270 31670 6310 31730
rect 2170 31660 6310 31670
rect 6380 31380 11240 31400
rect 6380 31320 6470 31380
rect 6530 31320 6580 31380
rect 6640 31320 6690 31380
rect 6750 31320 6800 31380
rect 6860 31320 6910 31380
rect 6970 31320 7020 31380
rect 7080 31320 7130 31380
rect 7190 31320 7240 31380
rect 7300 31320 7350 31380
rect 7410 31320 7460 31380
rect 7520 31320 7570 31380
rect 7630 31320 7680 31380
rect 7740 31320 7790 31380
rect 7850 31320 7900 31380
rect 7960 31320 8010 31380
rect 8070 31320 8120 31380
rect 8180 31320 8230 31380
rect 8290 31320 8340 31380
rect 8400 31320 8450 31380
rect 8510 31320 8560 31380
rect 8620 31320 8670 31380
rect 8730 31320 8780 31380
rect 8840 31320 8890 31380
rect 8950 31320 9000 31380
rect 9060 31320 9110 31380
rect 9170 31320 9220 31380
rect 9280 31320 9330 31380
rect 9390 31320 9440 31380
rect 9500 31320 9550 31380
rect 9610 31320 9660 31380
rect 9720 31320 9770 31380
rect 9830 31320 9880 31380
rect 9940 31320 9990 31380
rect 10050 31320 10100 31380
rect 10160 31320 10210 31380
rect 10270 31320 10320 31380
rect 10380 31320 10430 31380
rect 10490 31320 10540 31380
rect 10600 31320 10650 31380
rect 10710 31320 10760 31380
rect 10820 31320 10880 31380
rect 10940 31320 10990 31380
rect 11050 31320 11100 31380
rect 11160 31320 11240 31380
rect 6380 31300 11240 31320
rect 14830 30130 25680 30140
rect 14830 30060 14870 30130
rect 14930 30060 14970 30130
rect 15030 30060 15070 30130
rect 15130 30060 15170 30130
rect 15230 30060 15270 30130
rect 15330 30060 15370 30130
rect 15430 30060 15470 30130
rect 15530 30060 15570 30130
rect 15630 30060 15670 30130
rect 15730 30060 15780 30130
rect 15840 30060 15880 30130
rect 15940 30060 15990 30130
rect 16050 30060 16130 30130
rect 16190 30060 16270 30130
rect 16330 30060 16370 30130
rect 16430 30060 16470 30130
rect 16530 30060 16570 30130
rect 16630 30060 16670 30130
rect 16730 30060 16770 30130
rect 16830 30060 16870 30130
rect 16930 30060 16970 30130
rect 17030 30060 17070 30130
rect 17130 30060 17170 30130
rect 17230 30060 17270 30130
rect 17330 30060 17370 30130
rect 17430 30060 17470 30130
rect 17530 30060 17570 30130
rect 17630 30060 17670 30130
rect 17730 30060 17770 30130
rect 17830 30060 17870 30130
rect 17930 30060 17970 30130
rect 18030 30060 18070 30130
rect 18130 30060 18170 30130
rect 18230 30060 18270 30130
rect 18330 30060 18370 30130
rect 18430 30060 18470 30130
rect 18530 30060 18570 30130
rect 18630 30060 18670 30130
rect 18730 30060 18770 30130
rect 18830 30060 18870 30130
rect 18930 30060 18970 30130
rect 19030 30060 19070 30130
rect 19130 30060 19170 30130
rect 19230 30060 19270 30130
rect 19330 30060 19370 30130
rect 19430 30060 19470 30130
rect 19530 30060 19570 30130
rect 19630 30060 19670 30130
rect 19730 30060 19770 30130
rect 19830 30060 19870 30130
rect 19930 30060 19970 30130
rect 20030 30060 20070 30130
rect 20130 30060 20170 30130
rect 20230 30060 20270 30130
rect 20330 30060 20370 30130
rect 20430 30060 20470 30130
rect 20530 30060 20570 30130
rect 20630 30060 20670 30130
rect 20730 30060 20770 30130
rect 20830 30060 20870 30130
rect 20930 30060 20970 30130
rect 21030 30060 21070 30130
rect 21130 30060 21170 30130
rect 21230 30060 21270 30130
rect 21330 30060 21370 30130
rect 21430 30060 21470 30130
rect 21530 30060 21570 30130
rect 21630 30060 21670 30130
rect 21730 30060 21770 30130
rect 21830 30060 21870 30130
rect 21930 30060 21970 30130
rect 22030 30060 22070 30130
rect 22130 30060 22170 30130
rect 22230 30060 22270 30130
rect 22330 30060 22370 30130
rect 22430 30060 22470 30130
rect 22530 30060 22570 30130
rect 22630 30060 22670 30130
rect 22730 30060 22770 30130
rect 22830 30060 22870 30130
rect 22930 30060 22970 30130
rect 23030 30060 23070 30130
rect 23130 30060 23170 30130
rect 23230 30060 23270 30130
rect 23330 30060 23370 30130
rect 23430 30060 23470 30130
rect 23530 30060 23570 30130
rect 23630 30060 23670 30130
rect 23730 30060 23770 30130
rect 23830 30060 23870 30130
rect 23930 30060 23970 30130
rect 24030 30060 24070 30130
rect 24130 30060 24170 30130
rect 24230 30060 24270 30130
rect 24330 30060 24370 30130
rect 24430 30060 24470 30130
rect 24530 30060 24570 30130
rect 24630 30060 24670 30130
rect 24730 30060 24770 30130
rect 24830 30060 24870 30130
rect 24930 30060 24970 30130
rect 25030 30060 25070 30130
rect 25130 30060 25170 30130
rect 25230 30060 25270 30130
rect 25330 30060 25370 30130
rect 25430 30060 25470 30130
rect 25530 30060 25570 30130
rect 25630 30060 25680 30130
rect 14830 30050 25680 30060
rect 7280 24290 20620 24300
rect 7280 24250 7320 24290
rect 7360 24250 7400 24290
rect 7440 24250 7480 24290
rect 7520 24250 7560 24290
rect 7600 24250 7640 24290
rect 7680 24250 7720 24290
rect 7760 24250 7800 24290
rect 7840 24250 7890 24290
rect 7930 24250 7970 24290
rect 8010 24250 8050 24290
rect 8090 24250 8130 24290
rect 8170 24250 8210 24290
rect 8250 24250 8290 24290
rect 8330 24250 8400 24290
rect 8440 24250 8520 24290
rect 8560 24250 8600 24290
rect 8640 24250 8680 24290
rect 8720 24250 8760 24290
rect 8800 24250 8840 24290
rect 8880 24250 8920 24290
rect 8960 24250 9000 24290
rect 9040 24250 9080 24290
rect 9120 24250 9160 24290
rect 9200 24250 9270 24290
rect 9310 24250 9350 24290
rect 9390 24250 9430 24290
rect 9470 24250 9510 24290
rect 9550 24250 9590 24290
rect 9630 24250 9670 24290
rect 9710 24250 9750 24290
rect 9790 24250 9830 24290
rect 9870 24250 9910 24290
rect 9950 24250 9990 24290
rect 10030 24250 10070 24290
rect 10110 24250 10150 24290
rect 10190 24250 10230 24290
rect 10270 24250 10310 24290
rect 10350 24250 10390 24290
rect 10430 24250 10470 24290
rect 10510 24250 10550 24290
rect 10590 24250 10630 24290
rect 10670 24250 10710 24290
rect 10750 24250 10790 24290
rect 10830 24250 10870 24290
rect 10910 24250 10950 24290
rect 10990 24250 11030 24290
rect 11070 24250 11110 24290
rect 11150 24250 11190 24290
rect 11230 24250 11270 24290
rect 11310 24250 11350 24290
rect 11390 24250 11430 24290
rect 11470 24250 11510 24290
rect 11550 24250 11590 24290
rect 11630 24250 11670 24290
rect 11710 24250 11750 24290
rect 11790 24250 11830 24290
rect 11870 24250 11910 24290
rect 11950 24250 11990 24290
rect 12030 24250 12070 24290
rect 12110 24250 12150 24290
rect 12190 24250 12230 24290
rect 12270 24250 12310 24290
rect 12350 24250 12390 24290
rect 12430 24250 12470 24290
rect 12510 24250 12550 24290
rect 12590 24250 12630 24290
rect 12670 24250 12710 24290
rect 12750 24250 12790 24290
rect 12830 24250 12870 24290
rect 12910 24250 12950 24290
rect 12990 24250 13030 24290
rect 13070 24250 13110 24290
rect 13150 24250 13190 24290
rect 13230 24250 13270 24290
rect 13310 24250 13350 24290
rect 13390 24250 13430 24290
rect 13470 24250 13510 24290
rect 13550 24250 13590 24290
rect 13630 24250 13670 24290
rect 13710 24250 13750 24290
rect 13790 24250 13830 24290
rect 13870 24250 13910 24290
rect 13950 24250 13990 24290
rect 14030 24250 14070 24290
rect 14110 24250 14150 24290
rect 14190 24250 14230 24290
rect 14270 24250 14310 24290
rect 14350 24250 14390 24290
rect 14430 24250 14470 24290
rect 14510 24250 14550 24290
rect 14590 24250 14630 24290
rect 14670 24250 14710 24290
rect 14750 24250 14790 24290
rect 14830 24250 14870 24290
rect 14910 24250 14950 24290
rect 14990 24250 15030 24290
rect 15070 24250 15110 24290
rect 15150 24250 15190 24290
rect 15230 24250 15270 24290
rect 15310 24250 15350 24290
rect 15390 24250 15430 24290
rect 15470 24250 15510 24290
rect 15550 24250 15590 24290
rect 15630 24250 15670 24290
rect 15710 24250 15750 24290
rect 15790 24250 15830 24290
rect 15870 24250 15910 24290
rect 15950 24250 15990 24290
rect 16030 24250 16070 24290
rect 16110 24250 16150 24290
rect 16190 24250 16230 24290
rect 16270 24250 16310 24290
rect 16350 24250 16390 24290
rect 16430 24250 16470 24290
rect 16510 24250 16550 24290
rect 16590 24250 16630 24290
rect 16670 24250 16710 24290
rect 16750 24250 16790 24290
rect 16830 24250 16870 24290
rect 16910 24250 16950 24290
rect 16990 24250 17030 24290
rect 17070 24250 17110 24290
rect 17150 24250 17190 24290
rect 17230 24250 17270 24290
rect 17310 24250 17350 24290
rect 17390 24250 17430 24290
rect 17470 24250 17510 24290
rect 17550 24250 17590 24290
rect 17630 24250 17670 24290
rect 17710 24250 17750 24290
rect 17790 24250 17830 24290
rect 17870 24250 17910 24290
rect 17950 24250 17990 24290
rect 18030 24250 18070 24290
rect 18110 24250 18150 24290
rect 18190 24250 18230 24290
rect 18270 24250 18310 24290
rect 18350 24250 18390 24290
rect 18430 24250 18470 24290
rect 18510 24250 18550 24290
rect 18590 24250 18630 24290
rect 18670 24250 18710 24290
rect 18750 24250 18790 24290
rect 18830 24250 18870 24290
rect 18910 24250 18950 24290
rect 18990 24250 19030 24290
rect 19070 24250 19110 24290
rect 19150 24250 19190 24290
rect 19230 24250 19270 24290
rect 19310 24250 19350 24290
rect 19390 24250 19430 24290
rect 19470 24250 19510 24290
rect 19550 24250 19590 24290
rect 19630 24250 19670 24290
rect 19710 24250 19750 24290
rect 19790 24250 19830 24290
rect 19870 24250 19910 24290
rect 19950 24250 19990 24290
rect 20030 24250 20070 24290
rect 20110 24250 20150 24290
rect 20190 24250 20230 24290
rect 20270 24250 20310 24290
rect 20350 24250 20390 24290
rect 20430 24250 20470 24290
rect 20510 24250 20550 24290
rect 20590 24250 20620 24290
rect 7280 24240 20620 24250
rect 7280 23320 20620 23330
rect 7280 23280 7310 23320
rect 7350 23280 7390 23320
rect 7430 23280 7470 23320
rect 7510 23280 7550 23320
rect 7590 23280 7630 23320
rect 7670 23280 7710 23320
rect 7750 23280 7790 23320
rect 7830 23280 7870 23320
rect 7910 23280 7950 23320
rect 7990 23280 8030 23320
rect 8070 23280 8110 23320
rect 8150 23280 8190 23320
rect 8230 23280 8270 23320
rect 8310 23280 8350 23320
rect 8390 23280 8430 23320
rect 8470 23280 8520 23320
rect 8560 23280 8600 23320
rect 8640 23280 8680 23320
rect 8720 23280 8760 23320
rect 8800 23280 8840 23320
rect 8880 23280 8920 23320
rect 8960 23280 9000 23320
rect 9040 23280 9080 23320
rect 9120 23280 9160 23320
rect 9200 23280 9270 23320
rect 9310 23280 9350 23320
rect 9390 23280 9430 23320
rect 9470 23280 9510 23320
rect 9550 23280 9590 23320
rect 9630 23280 9670 23320
rect 9710 23280 9750 23320
rect 9790 23280 9830 23320
rect 9870 23280 9910 23320
rect 9950 23280 9990 23320
rect 10030 23280 10070 23320
rect 10110 23280 10150 23320
rect 10190 23280 10230 23320
rect 10270 23280 10310 23320
rect 10350 23280 10390 23320
rect 10430 23280 10470 23320
rect 10510 23280 10550 23320
rect 10590 23280 10630 23320
rect 10670 23280 10710 23320
rect 10750 23280 10790 23320
rect 10830 23280 10870 23320
rect 10910 23280 10950 23320
rect 10990 23280 11030 23320
rect 11070 23280 11110 23320
rect 11150 23280 11190 23320
rect 11230 23280 11270 23320
rect 11310 23280 11350 23320
rect 11390 23280 11430 23320
rect 11470 23280 11510 23320
rect 11550 23280 11590 23320
rect 11630 23280 11670 23320
rect 11710 23280 11750 23320
rect 11790 23280 11830 23320
rect 11870 23280 11910 23320
rect 11950 23280 11990 23320
rect 12030 23280 12070 23320
rect 12110 23280 12150 23320
rect 12190 23280 12230 23320
rect 12270 23280 12310 23320
rect 12350 23280 12390 23320
rect 12430 23280 12470 23320
rect 12510 23280 12550 23320
rect 12590 23280 12630 23320
rect 12670 23280 12710 23320
rect 12750 23280 12790 23320
rect 12830 23280 12870 23320
rect 12910 23280 12950 23320
rect 12990 23280 13030 23320
rect 13070 23280 13110 23320
rect 13150 23280 13190 23320
rect 13230 23280 13270 23320
rect 13310 23280 13350 23320
rect 13390 23280 13430 23320
rect 13470 23280 13510 23320
rect 13550 23280 13590 23320
rect 13630 23280 13670 23320
rect 13710 23280 13750 23320
rect 13790 23280 13830 23320
rect 13870 23280 13910 23320
rect 13950 23280 13990 23320
rect 14030 23280 14070 23320
rect 14110 23280 14150 23320
rect 14190 23280 14230 23320
rect 14270 23280 14310 23320
rect 14350 23280 14390 23320
rect 14430 23280 14470 23320
rect 14510 23280 14550 23320
rect 14590 23280 14630 23320
rect 14670 23280 14710 23320
rect 14750 23280 14790 23320
rect 14830 23280 14870 23320
rect 14910 23280 14950 23320
rect 14990 23280 15030 23320
rect 15070 23280 15110 23320
rect 15150 23280 15190 23320
rect 15230 23280 15270 23320
rect 15310 23280 15350 23320
rect 15390 23280 15430 23320
rect 15470 23280 15510 23320
rect 15550 23280 15590 23320
rect 15630 23280 15670 23320
rect 15710 23280 15750 23320
rect 15790 23280 15830 23320
rect 15870 23280 15910 23320
rect 15950 23280 15990 23320
rect 16030 23280 16070 23320
rect 16110 23280 16150 23320
rect 16190 23280 16230 23320
rect 16270 23280 16310 23320
rect 16350 23280 16390 23320
rect 16430 23280 16470 23320
rect 16510 23280 16550 23320
rect 16590 23280 16630 23320
rect 16670 23280 16710 23320
rect 16750 23280 16790 23320
rect 16830 23280 16870 23320
rect 16910 23280 16950 23320
rect 16990 23280 17030 23320
rect 17070 23280 17110 23320
rect 17150 23280 17190 23320
rect 17230 23280 17270 23320
rect 17310 23280 17350 23320
rect 17390 23280 17430 23320
rect 17470 23280 17510 23320
rect 17550 23280 17590 23320
rect 17630 23280 17670 23320
rect 17710 23280 17750 23320
rect 17790 23280 17830 23320
rect 17870 23280 17910 23320
rect 17950 23280 17990 23320
rect 18030 23280 18070 23320
rect 18110 23280 18150 23320
rect 18190 23280 18230 23320
rect 18270 23280 18310 23320
rect 18350 23280 18390 23320
rect 18430 23280 18470 23320
rect 18510 23280 18550 23320
rect 18590 23280 18630 23320
rect 18670 23280 18710 23320
rect 18750 23280 18790 23320
rect 18830 23280 18870 23320
rect 18910 23280 18950 23320
rect 18990 23280 19030 23320
rect 19070 23280 19110 23320
rect 19150 23280 19190 23320
rect 19230 23280 19270 23320
rect 19310 23280 19350 23320
rect 19390 23280 19430 23320
rect 19470 23280 19510 23320
rect 19550 23280 19590 23320
rect 19630 23280 19670 23320
rect 19710 23280 19750 23320
rect 19790 23280 19830 23320
rect 19870 23280 19910 23320
rect 19950 23280 19990 23320
rect 20030 23280 20070 23320
rect 20110 23280 20150 23320
rect 20190 23280 20230 23320
rect 20270 23280 20310 23320
rect 20350 23280 20390 23320
rect 20430 23280 20470 23320
rect 20510 23280 20550 23320
rect 20590 23280 20620 23320
rect 7280 23270 20620 23280
rect 7280 17700 20620 17710
rect 7280 17660 7320 17700
rect 7360 17660 7400 17700
rect 7440 17660 7480 17700
rect 7520 17660 7560 17700
rect 7600 17660 7640 17700
rect 7680 17660 7720 17700
rect 7760 17660 7800 17700
rect 7840 17660 7880 17700
rect 7920 17660 7960 17700
rect 8000 17660 8040 17700
rect 8080 17660 8120 17700
rect 8160 17660 8200 17700
rect 8240 17660 8280 17700
rect 8320 17660 8360 17700
rect 8400 17660 8440 17700
rect 8480 17660 8520 17700
rect 8560 17660 8600 17700
rect 8640 17660 8680 17700
rect 8720 17660 8760 17700
rect 8800 17660 8840 17700
rect 8880 17660 8920 17700
rect 8960 17660 9000 17700
rect 9040 17660 9080 17700
rect 9120 17660 9160 17700
rect 9200 17660 9270 17700
rect 9310 17660 9350 17700
rect 9390 17660 9430 17700
rect 9470 17660 9510 17700
rect 9550 17660 9590 17700
rect 9630 17660 9670 17700
rect 9710 17660 9750 17700
rect 9790 17660 9830 17700
rect 9870 17660 9910 17700
rect 9950 17660 9990 17700
rect 10030 17660 10070 17700
rect 10110 17660 10150 17700
rect 10190 17660 10230 17700
rect 10270 17660 10310 17700
rect 10350 17660 10390 17700
rect 10430 17660 10470 17700
rect 10510 17660 10550 17700
rect 10590 17660 10630 17700
rect 10670 17660 10710 17700
rect 10750 17660 10790 17700
rect 10830 17660 10870 17700
rect 10910 17660 10950 17700
rect 10990 17660 11030 17700
rect 11070 17660 11110 17700
rect 11150 17660 11190 17700
rect 11230 17660 11270 17700
rect 11310 17660 11350 17700
rect 11390 17660 11430 17700
rect 11470 17660 11510 17700
rect 11550 17660 11590 17700
rect 11630 17660 11670 17700
rect 11710 17660 11750 17700
rect 11790 17660 11830 17700
rect 11870 17660 11910 17700
rect 11950 17660 11990 17700
rect 12030 17660 12070 17700
rect 12110 17660 12150 17700
rect 12190 17660 12230 17700
rect 12270 17660 12310 17700
rect 12350 17660 12390 17700
rect 12430 17660 12470 17700
rect 12510 17660 12550 17700
rect 12590 17660 12630 17700
rect 12670 17660 12710 17700
rect 12750 17660 12790 17700
rect 12830 17660 12870 17700
rect 12910 17660 12950 17700
rect 12990 17660 13030 17700
rect 13070 17660 13110 17700
rect 13150 17660 13190 17700
rect 13230 17660 13270 17700
rect 13310 17660 13350 17700
rect 13390 17660 13430 17700
rect 13470 17660 13510 17700
rect 13550 17660 13590 17700
rect 13630 17660 13670 17700
rect 13710 17660 13750 17700
rect 13790 17660 13830 17700
rect 13870 17660 13910 17700
rect 13950 17660 13990 17700
rect 14030 17660 14070 17700
rect 14110 17660 14150 17700
rect 14190 17660 14230 17700
rect 14270 17660 14310 17700
rect 14350 17660 14390 17700
rect 14430 17660 14470 17700
rect 14510 17660 14550 17700
rect 14590 17660 14630 17700
rect 14670 17660 14710 17700
rect 14750 17660 14790 17700
rect 14830 17660 14870 17700
rect 14910 17660 14950 17700
rect 14990 17660 15030 17700
rect 15070 17660 15110 17700
rect 15150 17660 15190 17700
rect 15230 17660 15270 17700
rect 15310 17660 15350 17700
rect 15390 17660 15430 17700
rect 15470 17660 15510 17700
rect 15550 17660 15590 17700
rect 15630 17660 15670 17700
rect 15710 17660 15750 17700
rect 15790 17660 15830 17700
rect 15870 17660 15910 17700
rect 15950 17660 15990 17700
rect 16030 17660 16070 17700
rect 16110 17660 16150 17700
rect 16190 17660 16230 17700
rect 16270 17660 16310 17700
rect 16350 17660 16390 17700
rect 16430 17660 16470 17700
rect 16510 17660 16550 17700
rect 16590 17660 16630 17700
rect 16670 17660 16710 17700
rect 16750 17660 16790 17700
rect 16830 17660 16870 17700
rect 16910 17660 16950 17700
rect 16990 17660 17030 17700
rect 17070 17660 17110 17700
rect 17150 17660 17190 17700
rect 17230 17660 17270 17700
rect 17310 17660 17350 17700
rect 17390 17660 17430 17700
rect 17470 17660 17510 17700
rect 17550 17660 17590 17700
rect 17630 17660 17670 17700
rect 17710 17660 17750 17700
rect 17790 17660 17830 17700
rect 17870 17660 17910 17700
rect 17950 17660 17990 17700
rect 18030 17660 18070 17700
rect 18110 17660 18150 17700
rect 18190 17660 18230 17700
rect 18270 17660 18310 17700
rect 18350 17660 18390 17700
rect 18430 17660 18470 17700
rect 18510 17660 18550 17700
rect 18590 17660 18630 17700
rect 18670 17660 18710 17700
rect 18750 17660 18790 17700
rect 18830 17660 18870 17700
rect 18910 17660 18950 17700
rect 18990 17660 19030 17700
rect 19070 17660 19110 17700
rect 19150 17660 19190 17700
rect 19230 17660 19270 17700
rect 19310 17660 19350 17700
rect 19390 17660 19430 17700
rect 19470 17660 19510 17700
rect 19550 17660 19590 17700
rect 19630 17660 19670 17700
rect 19710 17660 19750 17700
rect 19790 17660 19830 17700
rect 19870 17660 19910 17700
rect 19950 17660 19990 17700
rect 20030 17660 20070 17700
rect 20110 17660 20150 17700
rect 20190 17660 20230 17700
rect 20270 17660 20310 17700
rect 20350 17660 20390 17700
rect 20430 17660 20470 17700
rect 20510 17660 20550 17700
rect 20590 17660 20620 17700
rect 7280 17650 20620 17660
rect 9620 15660 21160 15670
rect 9620 15620 9710 15660
rect 9750 15620 9790 15660
rect 9830 15620 9870 15660
rect 9910 15620 9950 15660
rect 9990 15620 10030 15660
rect 10070 15620 10110 15660
rect 10150 15620 10190 15660
rect 10230 15620 10270 15660
rect 10310 15620 10350 15660
rect 10390 15620 10430 15660
rect 10470 15620 10510 15660
rect 10550 15620 10590 15660
rect 10630 15620 10670 15660
rect 10710 15620 10750 15660
rect 10790 15620 10830 15660
rect 10870 15620 10910 15660
rect 10950 15620 10990 15660
rect 11030 15620 11070 15660
rect 11110 15620 11150 15660
rect 11190 15620 11230 15660
rect 11270 15620 11310 15660
rect 11350 15620 11390 15660
rect 11430 15620 11470 15660
rect 11510 15620 11550 15660
rect 11590 15620 11630 15660
rect 11670 15620 11710 15660
rect 11750 15620 11790 15660
rect 11830 15620 11870 15660
rect 11910 15620 11950 15660
rect 11990 15620 12030 15660
rect 12070 15620 12110 15660
rect 12150 15620 12190 15660
rect 12230 15620 12270 15660
rect 12310 15620 12350 15660
rect 12390 15620 12430 15660
rect 12470 15620 12510 15660
rect 12550 15620 12590 15660
rect 12630 15620 12670 15660
rect 12710 15620 12750 15660
rect 12790 15620 12830 15660
rect 12870 15620 12910 15660
rect 12950 15620 12990 15660
rect 13030 15620 13070 15660
rect 13110 15620 13150 15660
rect 13190 15620 13230 15660
rect 13270 15620 13310 15660
rect 13350 15620 13390 15660
rect 13430 15620 13470 15660
rect 13510 15620 13550 15660
rect 13590 15620 13630 15660
rect 13670 15620 13710 15660
rect 13750 15620 13790 15660
rect 13830 15620 13870 15660
rect 13910 15620 13950 15660
rect 13990 15620 14030 15660
rect 14070 15620 14110 15660
rect 14150 15620 14190 15660
rect 14230 15620 14270 15660
rect 14310 15620 14350 15660
rect 14390 15620 14430 15660
rect 14470 15620 14510 15660
rect 14550 15620 14590 15660
rect 14630 15620 14670 15660
rect 14710 15620 14750 15660
rect 14790 15620 14830 15660
rect 14870 15620 14910 15660
rect 14950 15620 14990 15660
rect 15030 15620 15070 15660
rect 15110 15620 15150 15660
rect 15190 15620 15230 15660
rect 15270 15620 15310 15660
rect 15350 15620 15390 15660
rect 15430 15620 15470 15660
rect 15510 15620 15550 15660
rect 15590 15620 15630 15660
rect 15670 15620 15710 15660
rect 15750 15620 15790 15660
rect 15830 15620 15870 15660
rect 15910 15620 15950 15660
rect 15990 15620 16030 15660
rect 16070 15620 16110 15660
rect 16150 15620 16190 15660
rect 16230 15620 16270 15660
rect 16310 15620 16350 15660
rect 16390 15620 16430 15660
rect 16470 15620 16510 15660
rect 16550 15620 16590 15660
rect 16630 15620 16670 15660
rect 16710 15620 16750 15660
rect 16790 15620 16830 15660
rect 16870 15620 16910 15660
rect 16950 15620 16990 15660
rect 17030 15620 17070 15660
rect 17110 15620 17150 15660
rect 17190 15620 17230 15660
rect 17270 15620 17310 15660
rect 17350 15620 17390 15660
rect 17430 15620 17470 15660
rect 17510 15620 17550 15660
rect 17590 15620 17630 15660
rect 17670 15620 17710 15660
rect 17750 15620 17790 15660
rect 17830 15620 17870 15660
rect 17910 15620 17950 15660
rect 17990 15620 18030 15660
rect 18070 15620 18110 15660
rect 18150 15620 18190 15660
rect 18230 15620 18270 15660
rect 18310 15620 18350 15660
rect 18390 15620 18430 15660
rect 18470 15620 18510 15660
rect 18550 15620 18590 15660
rect 18630 15620 18670 15660
rect 18710 15620 18750 15660
rect 18790 15620 18830 15660
rect 18870 15620 18910 15660
rect 18950 15620 18990 15660
rect 19030 15620 19070 15660
rect 19110 15620 19150 15660
rect 19190 15620 19230 15660
rect 19270 15620 19310 15660
rect 19350 15620 19390 15660
rect 19430 15620 19470 15660
rect 19510 15620 19550 15660
rect 19590 15620 19630 15660
rect 19670 15620 19710 15660
rect 19750 15620 19800 15660
rect 19840 15620 19880 15660
rect 19920 15620 19960 15660
rect 20000 15620 20040 15660
rect 20080 15620 20120 15660
rect 20160 15620 20200 15660
rect 20240 15620 20280 15660
rect 20320 15620 20370 15660
rect 20410 15620 20450 15660
rect 20490 15620 20530 15660
rect 20570 15620 20610 15660
rect 20650 15620 20690 15660
rect 20730 15620 20770 15660
rect 20810 15620 20850 15660
rect 20890 15620 20930 15660
rect 20970 15620 21010 15660
rect 21050 15620 21090 15660
rect 21130 15620 21160 15660
rect 9620 15610 21160 15620
rect 9730 12050 21160 12060
rect 9730 12010 9810 12050
rect 9850 12010 9890 12050
rect 9930 12010 9970 12050
rect 10010 12010 10050 12050
rect 10090 12010 10130 12050
rect 10170 12010 10210 12050
rect 10250 12010 10290 12050
rect 10330 12010 10370 12050
rect 10410 12010 10450 12050
rect 10490 12010 10530 12050
rect 10570 12010 10610 12050
rect 10650 12010 10690 12050
rect 10730 12010 10770 12050
rect 10810 12010 10850 12050
rect 10890 12010 10930 12050
rect 10970 12010 11010 12050
rect 11050 12010 11090 12050
rect 11130 12010 11170 12050
rect 11210 12010 11250 12050
rect 11290 12010 11330 12050
rect 11370 12010 11410 12050
rect 11450 12010 11490 12050
rect 11530 12010 11570 12050
rect 11610 12010 11650 12050
rect 11690 12010 11730 12050
rect 11770 12010 11810 12050
rect 11850 12010 11890 12050
rect 11930 12010 11970 12050
rect 12010 12010 12050 12050
rect 12090 12010 12130 12050
rect 12170 12010 12210 12050
rect 12250 12010 12290 12050
rect 12330 12010 12370 12050
rect 12410 12010 12450 12050
rect 12490 12010 12530 12050
rect 12570 12010 12610 12050
rect 12650 12010 12690 12050
rect 12730 12010 12770 12050
rect 12810 12010 12850 12050
rect 12890 12010 12930 12050
rect 12970 12010 13010 12050
rect 13050 12010 13090 12050
rect 13130 12010 13170 12050
rect 13210 12010 13250 12050
rect 13290 12010 13330 12050
rect 13440 12010 13480 12050
rect 13520 12010 13560 12050
rect 13600 12010 13640 12050
rect 13680 12010 13720 12050
rect 13760 12010 13800 12050
rect 13840 12010 13880 12050
rect 13920 12010 13960 12050
rect 14000 12010 14040 12050
rect 14080 12010 14120 12050
rect 14160 12010 14200 12050
rect 14240 12010 14280 12050
rect 14320 12010 14360 12050
rect 14400 12010 14440 12050
rect 14480 12010 14520 12050
rect 14560 12010 14600 12050
rect 14640 12010 14680 12050
rect 14720 12010 14760 12050
rect 14800 12010 14840 12050
rect 14880 12010 14920 12050
rect 14960 12010 15000 12050
rect 15040 12010 15080 12050
rect 15120 12010 15160 12050
rect 15200 12010 15240 12050
rect 15280 12010 15320 12050
rect 15360 12010 15400 12050
rect 15440 12010 15480 12050
rect 15520 12010 15560 12050
rect 15600 12010 15640 12050
rect 15680 12010 15720 12050
rect 15760 12010 15800 12050
rect 15840 12010 15880 12050
rect 15920 12010 15960 12050
rect 16000 12010 16040 12050
rect 16080 12010 16120 12050
rect 16160 12010 16200 12050
rect 16240 12010 16280 12050
rect 16320 12010 16360 12050
rect 16400 12010 16440 12050
rect 16480 12010 16520 12050
rect 16560 12010 16600 12050
rect 16640 12010 16680 12050
rect 16720 12010 16760 12050
rect 16800 12010 16840 12050
rect 16880 12010 16920 12050
rect 16960 12010 17000 12050
rect 17040 12010 17080 12050
rect 17120 12010 17160 12050
rect 17200 12010 17240 12050
rect 17280 12010 17320 12050
rect 17360 12010 17400 12050
rect 17440 12010 17480 12050
rect 17520 12010 17560 12050
rect 17600 12010 17640 12050
rect 17680 12010 17720 12050
rect 17760 12010 17800 12050
rect 17840 12010 17880 12050
rect 17920 12010 17960 12050
rect 18000 12010 18040 12050
rect 18080 12010 18120 12050
rect 18160 12010 18200 12050
rect 18240 12010 18280 12050
rect 18320 12010 18360 12050
rect 18400 12010 18440 12050
rect 18480 12010 18520 12050
rect 18560 12010 18600 12050
rect 18640 12010 18680 12050
rect 18720 12010 18760 12050
rect 18800 12010 18840 12050
rect 18880 12010 18920 12050
rect 18960 12010 19000 12050
rect 19040 12010 19080 12050
rect 19120 12010 19160 12050
rect 19200 12010 19240 12050
rect 19280 12010 19320 12050
rect 19360 12010 19400 12050
rect 19440 12010 19480 12050
rect 19520 12010 19560 12050
rect 19600 12010 19640 12050
rect 19680 12010 19720 12050
rect 19760 12010 19800 12050
rect 19840 12010 19890 12050
rect 19930 12010 19970 12050
rect 20010 12010 20050 12050
rect 20090 12010 20130 12050
rect 20170 12010 20210 12050
rect 20250 12010 20290 12050
rect 20330 12010 20370 12050
rect 20410 12010 20460 12050
rect 20500 12010 20540 12050
rect 20580 12010 20620 12050
rect 20660 12010 20700 12050
rect 20740 12010 20780 12050
rect 20820 12010 20860 12050
rect 20900 12010 20940 12050
rect 20980 12010 21020 12050
rect 21060 12010 21160 12050
rect 7280 12000 21160 12010
rect 7280 11960 7330 12000
rect 7370 11960 7410 12000
rect 7450 11960 7490 12000
rect 7530 11960 7570 12000
rect 7610 11960 7650 12000
rect 7690 11960 7730 12000
rect 7770 11960 7810 12000
rect 7850 11960 7890 12000
rect 7930 11960 7970 12000
rect 8010 11960 8050 12000
rect 8090 11960 8130 12000
rect 8170 11960 8210 12000
rect 8250 11960 8290 12000
rect 8330 11960 8370 12000
rect 8410 11960 8450 12000
rect 8490 11960 8530 12000
rect 8570 11960 8610 12000
rect 8650 11960 8690 12000
rect 8730 11960 8770 12000
rect 8810 11960 8850 12000
rect 8890 11960 8930 12000
rect 8970 11960 9010 12000
rect 9050 11960 9090 12000
rect 9130 11960 9170 12000
rect 9210 11960 9250 12000
rect 9290 11960 9330 12000
rect 9370 11960 9410 12000
rect 9450 11960 9490 12000
rect 9530 11960 9570 12000
rect 9610 11960 9650 12000
rect 9690 11960 9730 12000
rect 9770 11960 9800 12000
rect 7280 11950 9800 11960
rect 7660 11410 8600 11420
rect 7660 11370 7720 11410
rect 7760 11370 7800 11410
rect 7840 11370 7880 11410
rect 7920 11370 7960 11410
rect 8000 11370 8040 11410
rect 8080 11370 8120 11410
rect 8160 11370 8200 11410
rect 8240 11370 8280 11410
rect 8320 11370 8360 11410
rect 8400 11370 8440 11410
rect 8480 11370 8520 11410
rect 8560 11370 8600 11410
rect 7660 11360 8600 11370
rect 7660 11330 7720 11360
rect 7660 11290 7670 11330
rect 7710 11290 7720 11330
rect 8540 11330 8600 11360
rect 7660 11250 7720 11290
rect 7660 11210 7670 11250
rect 7710 11210 7720 11250
rect 7660 11170 7720 11210
rect 7660 11130 7670 11170
rect 7710 11130 7720 11170
rect 7660 11100 7720 11130
rect 8540 11290 8550 11330
rect 8590 11290 8600 11330
rect 8540 11250 8600 11290
rect 8540 11210 8550 11250
rect 8590 11210 8600 11250
rect 8540 11170 8600 11210
rect 8540 11130 8550 11170
rect 8590 11130 8600 11170
rect 8540 11100 8600 11130
rect 7280 11090 7720 11100
rect 7280 11050 7330 11090
rect 7370 11050 7410 11090
rect 7450 11050 7490 11090
rect 7530 11050 7570 11090
rect 7610 11050 7650 11090
rect 7690 11050 7720 11090
rect 7280 11040 7720 11050
rect 8540 11090 9800 11100
rect 8540 11050 8610 11090
rect 8650 11050 8690 11090
rect 8730 11050 8770 11090
rect 8810 11050 8850 11090
rect 8890 11050 8930 11090
rect 8970 11050 9010 11090
rect 9050 11050 9090 11090
rect 9130 11050 9170 11090
rect 9210 11050 9250 11090
rect 9290 11050 9330 11090
rect 9370 11050 9410 11090
rect 9450 11050 9490 11090
rect 9530 11050 9570 11090
rect 9610 11050 9650 11090
rect 9690 11050 9730 11090
rect 9770 11050 9800 11090
rect 8540 11040 21160 11050
rect 9730 11000 9810 11040
rect 9850 11000 9890 11040
rect 9930 11000 9970 11040
rect 10010 11000 10050 11040
rect 10090 11000 10130 11040
rect 10170 11000 10210 11040
rect 10250 11000 10290 11040
rect 10330 11000 10370 11040
rect 10410 11000 10450 11040
rect 10490 11000 10530 11040
rect 10570 11000 10610 11040
rect 10650 11000 10690 11040
rect 10730 11000 10770 11040
rect 10810 11000 10850 11040
rect 10890 11000 10930 11040
rect 10970 11000 11010 11040
rect 11050 11000 11090 11040
rect 11130 11000 11170 11040
rect 11210 11000 11250 11040
rect 11290 11000 11330 11040
rect 11370 11000 11410 11040
rect 11450 11000 11490 11040
rect 11530 11000 11570 11040
rect 11610 11000 11650 11040
rect 11690 11000 11730 11040
rect 11770 11000 11810 11040
rect 11850 11000 11890 11040
rect 11930 11000 11970 11040
rect 12010 11000 12050 11040
rect 12090 11000 12130 11040
rect 12170 11000 12210 11040
rect 12250 11000 12290 11040
rect 12330 11000 12370 11040
rect 12410 11000 12450 11040
rect 12490 11000 12530 11040
rect 12570 11000 12610 11040
rect 12650 11000 12690 11040
rect 12730 11000 12770 11040
rect 12810 11000 12850 11040
rect 12890 11000 12930 11040
rect 12970 11000 13010 11040
rect 13050 11000 13090 11040
rect 13130 11000 13170 11040
rect 13210 11000 13250 11040
rect 13290 11000 13330 11040
rect 13410 11000 13450 11040
rect 13490 11000 13530 11040
rect 13570 11000 13610 11040
rect 13650 11000 13690 11040
rect 13730 11000 13770 11040
rect 13810 11000 13850 11040
rect 13890 11000 13930 11040
rect 13970 11000 14010 11040
rect 14050 11000 14090 11040
rect 14130 11000 14170 11040
rect 14210 11000 14250 11040
rect 14290 11000 14330 11040
rect 14370 11000 14410 11040
rect 14450 11000 14490 11040
rect 14530 11000 14570 11040
rect 14610 11000 14650 11040
rect 14690 11000 14730 11040
rect 14770 11000 14810 11040
rect 14850 11000 14890 11040
rect 14930 11000 14970 11040
rect 15010 11000 15050 11040
rect 15090 11000 15130 11040
rect 15170 11000 15210 11040
rect 15250 11000 15290 11040
rect 15330 11000 15370 11040
rect 15410 11000 15450 11040
rect 15490 11000 15530 11040
rect 15570 11000 15610 11040
rect 15650 11000 15690 11040
rect 15730 11000 15770 11040
rect 15810 11000 15850 11040
rect 15890 11000 15930 11040
rect 15970 11000 16010 11040
rect 16050 11000 16090 11040
rect 16130 11000 16170 11040
rect 16210 11000 16250 11040
rect 16290 11000 16330 11040
rect 16370 11000 16410 11040
rect 16450 11000 16490 11040
rect 16530 11000 16570 11040
rect 16610 11000 16650 11040
rect 16690 11000 16730 11040
rect 16770 11000 16810 11040
rect 16850 11000 16890 11040
rect 16930 11000 16970 11040
rect 17010 11000 17050 11040
rect 17090 11000 17130 11040
rect 17170 11000 17210 11040
rect 17250 11000 17290 11040
rect 17330 11000 17370 11040
rect 17410 11000 17450 11040
rect 17490 11000 17530 11040
rect 17570 11000 17610 11040
rect 17650 11000 17690 11040
rect 17730 11000 17770 11040
rect 17810 11000 17850 11040
rect 17890 11000 17930 11040
rect 17970 11000 18010 11040
rect 18050 11000 18090 11040
rect 18130 11000 18170 11040
rect 18210 11000 18250 11040
rect 18290 11000 18330 11040
rect 18370 11000 18410 11040
rect 18450 11000 18490 11040
rect 18530 11000 18570 11040
rect 18610 11000 18650 11040
rect 18690 11000 18730 11040
rect 18770 11000 18810 11040
rect 18850 11000 18890 11040
rect 18930 11000 18970 11040
rect 19010 11000 19050 11040
rect 19090 11000 19130 11040
rect 19170 11000 19210 11040
rect 19250 11000 19290 11040
rect 19330 11000 19370 11040
rect 19410 11000 19450 11040
rect 19490 11000 19540 11040
rect 19580 11000 19620 11040
rect 19660 11000 19700 11040
rect 19740 11000 19780 11040
rect 19820 11000 19860 11040
rect 19900 11000 19940 11040
rect 19980 11000 20020 11040
rect 20060 11000 20110 11040
rect 20150 11000 20190 11040
rect 20230 11000 20270 11040
rect 20310 11000 20350 11040
rect 20390 11000 20430 11040
rect 20470 11000 20510 11040
rect 20550 11000 20590 11040
rect 20630 11000 20670 11040
rect 20710 11000 20750 11040
rect 20790 11000 20830 11040
rect 20870 11000 20910 11040
rect 20950 11000 20990 11040
rect 21030 11000 21070 11040
rect 21110 11000 21160 11040
rect 9730 10990 21160 11000
rect 13600 3000 17020 3010
rect 13600 2950 13630 3000
rect 13690 2950 13850 3000
rect 13910 2950 14070 3000
rect 14130 2950 14290 3000
rect 14350 2950 14510 3000
rect 14570 2950 14730 3000
rect 14790 2950 14950 3000
rect 15010 2950 15170 3000
rect 15230 2950 15390 3000
rect 15450 2950 15610 3000
rect 15670 2950 15830 3000
rect 15890 2950 16050 3000
rect 16110 2950 16270 3000
rect 16330 2950 16490 3000
rect 16550 2950 16710 3000
rect 16770 2950 17020 3000
rect 13600 2940 17020 2950
rect 24210 2720 24290 2770
rect 24210 2660 24220 2720
rect 24280 2660 24290 2720
rect 24210 2620 24290 2660
rect 24210 2560 24220 2620
rect 24280 2560 24290 2620
rect 24210 2520 24290 2560
rect 24210 2460 24220 2520
rect 24280 2460 24290 2520
rect 24210 2420 24290 2460
rect 24210 2360 24220 2420
rect 24280 2360 24290 2420
rect 24210 2320 24290 2360
rect 24210 2260 24220 2320
rect 24280 2260 24290 2320
rect 24210 2220 24290 2260
rect 24210 2160 24220 2220
rect 24280 2160 24290 2220
rect 24210 2120 24290 2160
rect 24210 2060 24220 2120
rect 24280 2060 24290 2120
rect 24210 2030 24290 2060
rect 9850 1920 17020 1930
rect 9850 1870 9890 1920
rect 9950 1870 10110 1920
rect 10170 1870 10330 1920
rect 10390 1870 10550 1920
rect 10610 1870 10770 1920
rect 10830 1870 10990 1920
rect 11050 1870 11210 1920
rect 11270 1870 11430 1920
rect 11490 1870 11650 1920
rect 11710 1870 11870 1920
rect 11930 1870 12090 1920
rect 12150 1870 12310 1920
rect 12370 1870 12530 1920
rect 12590 1870 12750 1920
rect 12810 1870 12970 1920
rect 13030 1870 13630 1920
rect 13690 1870 13850 1920
rect 13910 1870 14070 1920
rect 14130 1870 14290 1920
rect 14350 1870 14510 1920
rect 14570 1870 14730 1920
rect 14790 1870 14950 1920
rect 15010 1870 15170 1920
rect 15230 1870 15390 1920
rect 15450 1870 15610 1920
rect 15670 1870 15830 1920
rect 15890 1870 16050 1920
rect 16110 1870 16270 1920
rect 16330 1870 16490 1920
rect 16550 1870 16710 1920
rect 16770 1870 17020 1920
rect 9850 1860 17020 1870
<< nsubdiff >>
rect 21790 43350 23630 43360
rect 21790 43280 21830 43350
rect 21890 43280 21930 43350
rect 21990 43280 22030 43350
rect 22090 43280 22130 43350
rect 22190 43280 22230 43350
rect 22290 43280 22330 43350
rect 22390 43280 22430 43350
rect 22490 43280 22530 43350
rect 22590 43280 22630 43350
rect 22690 43280 22730 43350
rect 22790 43280 22830 43350
rect 22890 43280 22930 43350
rect 22990 43280 23030 43350
rect 23090 43280 23130 43350
rect 23190 43280 23230 43350
rect 23290 43280 23330 43350
rect 23390 43280 23430 43350
rect 23490 43280 23530 43350
rect 23590 43280 23630 43350
rect 21790 43270 23630 43280
rect 2439 42160 2999 42170
rect 2439 42110 2469 42160
rect 2519 42110 2559 42160
rect 2609 42110 2649 42160
rect 2699 42110 2739 42160
rect 2789 42110 2829 42160
rect 2879 42110 2919 42160
rect 2969 42110 2999 42160
rect 2439 42100 2999 42110
rect 5949 41970 9979 41980
rect 3390 41950 4329 41960
rect 3390 41900 3429 41950
rect 3479 41900 3519 41950
rect 3569 41900 3609 41950
rect 3659 41900 3699 41950
rect 3749 41900 3789 41950
rect 3839 41900 3879 41950
rect 3929 41900 3969 41950
rect 4019 41900 4059 41950
rect 4109 41900 4149 41950
rect 4199 41900 4239 41950
rect 4289 41900 4329 41950
rect 3390 41890 4329 41900
rect 4539 41950 5479 41960
rect 4539 41890 4579 41950
rect 4639 41890 5479 41950
rect 5949 41910 6009 41970
rect 6069 41910 6119 41970
rect 6179 41910 6229 41970
rect 6289 41910 6339 41970
rect 6399 41910 6449 41970
rect 6509 41910 6559 41970
rect 6619 41910 6669 41970
rect 6729 41910 6779 41970
rect 6839 41910 6889 41970
rect 6949 41910 6999 41970
rect 7059 41910 7109 41970
rect 7169 41910 7219 41970
rect 7279 41910 7329 41970
rect 7389 41910 7439 41970
rect 7499 41910 7549 41970
rect 7609 41910 7659 41970
rect 7719 41910 7769 41970
rect 7829 41910 7879 41970
rect 7939 41910 7989 41970
rect 8049 41910 8099 41970
rect 8159 41910 8209 41970
rect 8269 41910 8319 41970
rect 8379 41910 8429 41970
rect 8489 41910 8539 41970
rect 8599 41910 8649 41970
rect 8709 41910 8759 41970
rect 8819 41910 8869 41970
rect 8929 41910 8979 41970
rect 9039 41910 9089 41970
rect 9149 41910 9199 41970
rect 9259 41910 9309 41970
rect 9369 41910 9419 41970
rect 9479 41910 9529 41970
rect 9589 41910 9639 41970
rect 9699 41910 9749 41970
rect 9809 41910 9859 41970
rect 9919 41910 9979 41970
rect 5949 41900 9979 41910
rect 4539 41880 5479 41890
rect 3260 40670 4200 40680
rect 3260 40610 3320 40670
rect 3380 40610 3430 40670
rect 3490 40610 3540 40670
rect 3600 40610 3650 40670
rect 3710 40610 3760 40670
rect 3820 40610 3870 40670
rect 3930 40610 3980 40670
rect 4040 40610 4090 40670
rect 4150 40610 4200 40670
rect 3260 40600 4200 40610
rect 4539 40660 5429 40680
rect 4539 40620 4659 40660
rect 5399 40620 5429 40660
rect 4539 40600 5429 40620
rect 6349 40650 9969 40660
rect 6349 40590 6409 40650
rect 6469 40590 6519 40650
rect 6579 40590 6629 40650
rect 6689 40590 6739 40650
rect 6799 40590 6849 40650
rect 6909 40590 6959 40650
rect 7019 40590 7069 40650
rect 7129 40590 7179 40650
rect 7239 40590 7289 40650
rect 7349 40590 7399 40650
rect 7459 40590 7509 40650
rect 7569 40590 7619 40650
rect 7679 40590 7729 40650
rect 7789 40590 7839 40650
rect 7899 40590 7949 40650
rect 8009 40590 8059 40650
rect 8119 40590 8169 40650
rect 8229 40590 8279 40650
rect 8339 40590 8389 40650
rect 8449 40590 8499 40650
rect 8559 40590 8609 40650
rect 8669 40590 8719 40650
rect 8779 40590 8829 40650
rect 8889 40590 8939 40650
rect 8999 40590 9049 40650
rect 9109 40590 9159 40650
rect 9219 40590 9269 40650
rect 9329 40590 9379 40650
rect 9439 40590 9489 40650
rect 9549 40590 9599 40650
rect 9659 40590 9709 40650
rect 9769 40590 9819 40650
rect 9879 40590 9969 40650
rect 6349 40580 9969 40590
rect 15180 36340 24910 36350
rect 15180 36270 15220 36340
rect 15280 36270 15320 36340
rect 15380 36270 15420 36340
rect 15480 36270 15520 36340
rect 15580 36270 15620 36340
rect 15680 36270 15720 36340
rect 15780 36270 15820 36340
rect 15880 36270 15920 36340
rect 15980 36270 16020 36340
rect 16080 36270 16120 36340
rect 16180 36270 16220 36340
rect 16280 36270 16320 36340
rect 16380 36270 16420 36340
rect 16480 36270 16520 36340
rect 16580 36270 16620 36340
rect 16680 36270 16720 36340
rect 16780 36270 16820 36340
rect 16880 36270 16920 36340
rect 16980 36270 17020 36340
rect 17080 36270 17120 36340
rect 17180 36270 17220 36340
rect 17280 36270 17320 36340
rect 17380 36270 17420 36340
rect 17480 36270 17520 36340
rect 17580 36270 17620 36340
rect 17680 36270 17720 36340
rect 17780 36270 17820 36340
rect 17880 36270 17920 36340
rect 17980 36270 18020 36340
rect 18080 36270 18120 36340
rect 18180 36270 18220 36340
rect 18280 36270 18320 36340
rect 18380 36270 18420 36340
rect 18480 36270 18520 36340
rect 18580 36270 18620 36340
rect 18680 36270 18720 36340
rect 18780 36270 18820 36340
rect 18880 36270 18920 36340
rect 18980 36270 19020 36340
rect 19080 36270 19120 36340
rect 19180 36270 19220 36340
rect 19280 36270 19320 36340
rect 19380 36270 19420 36340
rect 19480 36270 19520 36340
rect 19580 36270 19620 36340
rect 19680 36270 19720 36340
rect 19780 36270 19820 36340
rect 19880 36270 19920 36340
rect 19980 36270 20020 36340
rect 20080 36270 20120 36340
rect 20180 36270 20220 36340
rect 20280 36270 20320 36340
rect 20380 36270 20420 36340
rect 20480 36270 20520 36340
rect 20580 36270 20620 36340
rect 20680 36270 20720 36340
rect 20780 36270 20820 36340
rect 20880 36270 20920 36340
rect 20980 36270 21020 36340
rect 21080 36270 21120 36340
rect 21180 36270 21220 36340
rect 21280 36270 21320 36340
rect 21380 36270 21420 36340
rect 21480 36270 21520 36340
rect 21580 36270 21620 36340
rect 21680 36270 21720 36340
rect 21780 36270 21820 36340
rect 21880 36270 21920 36340
rect 21980 36270 22020 36340
rect 22080 36270 22120 36340
rect 22180 36270 22220 36340
rect 22280 36270 22320 36340
rect 22380 36270 22420 36340
rect 22480 36270 22520 36340
rect 22580 36270 22620 36340
rect 22680 36270 22720 36340
rect 22780 36270 22820 36340
rect 22880 36270 22920 36340
rect 22980 36270 23020 36340
rect 23080 36270 23120 36340
rect 23180 36270 23220 36340
rect 23280 36270 23320 36340
rect 23380 36270 23420 36340
rect 23480 36270 23520 36340
rect 23580 36270 23620 36340
rect 23680 36270 23720 36340
rect 23780 36270 23820 36340
rect 23880 36270 23920 36340
rect 23980 36270 24020 36340
rect 24080 36270 24120 36340
rect 24180 36270 24220 36340
rect 24280 36270 24320 36340
rect 24380 36270 24420 36340
rect 24480 36270 24520 36340
rect 24580 36270 24620 36340
rect 24680 36270 24720 36340
rect 24780 36270 24820 36340
rect 24880 36270 24910 36340
rect 15180 36260 24910 36270
rect 15160 36110 15340 36120
rect 15160 36050 15200 36110
rect 15300 36050 15340 36110
rect 15160 36040 15340 36050
rect 6340 34040 10880 34050
rect 6340 33980 6380 34040
rect 6440 33980 6480 34040
rect 6540 33980 6580 34040
rect 6640 33980 6680 34040
rect 6740 33980 6780 34040
rect 6840 33980 6880 34040
rect 6940 33980 6980 34040
rect 7040 33980 7080 34040
rect 7140 33980 7180 34040
rect 7240 33980 7280 34040
rect 7340 33980 7380 34040
rect 7440 33980 7480 34040
rect 7540 33980 7580 34040
rect 7640 33980 7680 34040
rect 7740 33980 7780 34040
rect 7840 33980 7880 34040
rect 7940 33980 7980 34040
rect 8040 33980 8080 34040
rect 8140 33980 8180 34040
rect 8240 33980 8280 34040
rect 8340 33980 8380 34040
rect 8440 33980 8480 34040
rect 8540 33980 8580 34040
rect 8640 33980 8680 34040
rect 8740 33980 8780 34040
rect 8840 33980 8880 34040
rect 8940 33980 8980 34040
rect 9040 33980 9080 34040
rect 9140 33980 9180 34040
rect 9240 33980 9280 34040
rect 9340 33980 9380 34040
rect 9440 33980 9480 34040
rect 9540 33980 9580 34040
rect 9640 33980 9680 34040
rect 9740 33980 9780 34040
rect 9840 33980 9880 34040
rect 9940 33980 9980 34040
rect 10040 33980 10080 34040
rect 10140 33980 10180 34040
rect 10240 33980 10280 34040
rect 10340 33980 10380 34040
rect 10440 33980 10480 34040
rect 10540 33980 10580 34040
rect 10640 33980 10680 34040
rect 10740 33980 10780 34040
rect 10840 33980 10880 34040
rect 6340 33970 10880 33980
rect 3770 33620 6210 33630
rect 3770 33560 3810 33620
rect 3870 33560 3910 33620
rect 3970 33560 4010 33620
rect 4070 33560 4110 33620
rect 4170 33560 4210 33620
rect 4270 33560 4310 33620
rect 4370 33560 4410 33620
rect 4470 33560 4510 33620
rect 4570 33560 4610 33620
rect 4670 33560 4710 33620
rect 4770 33560 4810 33620
rect 4870 33560 4910 33620
rect 4970 33560 5010 33620
rect 5070 33560 5110 33620
rect 5170 33560 5210 33620
rect 5270 33560 5310 33620
rect 5370 33560 5410 33620
rect 5470 33560 5510 33620
rect 5570 33560 5610 33620
rect 5670 33560 5710 33620
rect 5770 33560 5810 33620
rect 5870 33560 5910 33620
rect 5970 33560 6010 33620
rect 6070 33560 6110 33620
rect 6170 33560 6210 33620
rect 3770 33550 6210 33560
rect 13728 32460 13888 32480
rect 13728 32420 13768 32460
rect 13848 32420 13888 32460
rect 13728 32400 13888 32420
rect 16030 32180 25410 32190
rect 16030 32110 16120 32180
rect 16180 32110 16220 32180
rect 16280 32110 16320 32180
rect 16380 32110 16420 32180
rect 16480 32110 16520 32180
rect 16580 32110 16620 32180
rect 16680 32110 16720 32180
rect 16780 32110 16820 32180
rect 16880 32110 16920 32180
rect 16980 32110 17020 32180
rect 17080 32110 17120 32180
rect 17180 32110 17220 32180
rect 17280 32110 17320 32180
rect 17380 32110 17420 32180
rect 17480 32110 17520 32180
rect 17580 32110 17620 32180
rect 17680 32110 17720 32180
rect 17780 32110 17820 32180
rect 17880 32110 17920 32180
rect 17980 32110 18020 32180
rect 18080 32110 18120 32180
rect 18180 32110 18220 32180
rect 18280 32110 18320 32180
rect 18380 32110 18420 32180
rect 18480 32110 18520 32180
rect 18580 32110 18620 32180
rect 18680 32110 18720 32180
rect 18780 32110 18820 32180
rect 18880 32110 18920 32180
rect 18980 32110 19020 32180
rect 19080 32110 19120 32180
rect 19180 32110 19220 32180
rect 19280 32110 19320 32180
rect 19380 32110 19420 32180
rect 19480 32110 19520 32180
rect 19580 32110 19620 32180
rect 19680 32110 19720 32180
rect 19780 32110 19820 32180
rect 19880 32110 19920 32180
rect 19980 32110 20020 32180
rect 20080 32110 20120 32180
rect 20180 32110 20220 32180
rect 20280 32110 20320 32180
rect 20380 32110 20420 32180
rect 20480 32110 20520 32180
rect 20580 32110 20620 32180
rect 20680 32110 20720 32180
rect 20780 32110 20820 32180
rect 20880 32110 20920 32180
rect 20980 32110 21020 32180
rect 21080 32110 21120 32180
rect 21180 32110 21220 32180
rect 21280 32110 21320 32180
rect 21380 32110 21420 32180
rect 21480 32110 21520 32180
rect 21580 32110 21620 32180
rect 21680 32110 21720 32180
rect 21780 32110 21820 32180
rect 21880 32110 21920 32180
rect 21980 32110 22020 32180
rect 22080 32110 22120 32180
rect 22180 32110 22220 32180
rect 22280 32110 22320 32180
rect 22380 32110 22420 32180
rect 22480 32110 22520 32180
rect 22580 32110 22620 32180
rect 22680 32110 22720 32180
rect 22780 32110 22820 32180
rect 22880 32110 22920 32180
rect 22980 32110 23020 32180
rect 23080 32110 23120 32180
rect 23180 32110 23220 32180
rect 23280 32110 23320 32180
rect 23380 32110 23420 32180
rect 23480 32110 23520 32180
rect 23580 32110 23620 32180
rect 23680 32110 23720 32180
rect 23780 32110 23820 32180
rect 23880 32110 23920 32180
rect 23980 32110 24020 32180
rect 24080 32110 24120 32180
rect 24180 32110 24220 32180
rect 24280 32110 24320 32180
rect 24380 32110 24420 32180
rect 24480 32110 24520 32180
rect 24580 32110 24620 32180
rect 24680 32110 24720 32180
rect 24780 32110 24820 32180
rect 24880 32110 24920 32180
rect 24980 32110 25020 32180
rect 25080 32110 25120 32180
rect 25180 32110 25220 32180
rect 25280 32110 25320 32180
rect 25380 32110 25410 32180
rect 16030 32100 25410 32110
rect 6400 29900 11240 29910
rect 6400 29840 6440 29900
rect 6500 29840 6540 29900
rect 6600 29840 6640 29900
rect 6700 29840 6740 29900
rect 6800 29840 6840 29900
rect 6900 29840 6940 29900
rect 7000 29840 7040 29900
rect 7100 29840 7140 29900
rect 7200 29840 7240 29900
rect 7300 29840 7340 29900
rect 7400 29840 7440 29900
rect 7500 29840 7540 29900
rect 7600 29840 7640 29900
rect 7700 29840 7740 29900
rect 7800 29840 7840 29900
rect 7900 29840 7940 29900
rect 8000 29840 8040 29900
rect 8100 29840 8140 29900
rect 8200 29840 8240 29900
rect 8300 29840 8340 29900
rect 8400 29840 8440 29900
rect 8500 29840 8540 29900
rect 8600 29840 8640 29900
rect 8700 29840 8740 29900
rect 8800 29840 8840 29900
rect 8900 29840 8940 29900
rect 9000 29840 9040 29900
rect 9100 29840 9140 29900
rect 9200 29840 9240 29900
rect 9300 29840 9340 29900
rect 9400 29840 9440 29900
rect 9500 29840 9540 29900
rect 9600 29840 9640 29900
rect 9700 29840 9740 29900
rect 9800 29840 9840 29900
rect 9900 29840 9940 29900
rect 10000 29840 10040 29900
rect 10100 29840 10140 29900
rect 10200 29840 10240 29900
rect 10300 29840 10340 29900
rect 10400 29840 10440 29900
rect 10500 29840 10540 29900
rect 10600 29840 10640 29900
rect 10700 29840 10740 29900
rect 10800 29840 10840 29900
rect 10900 29840 10940 29900
rect 11000 29840 11040 29900
rect 11100 29840 11140 29900
rect 11200 29840 11240 29900
rect 6400 29830 11240 29840
rect 2170 29370 6310 29380
rect 2170 29310 2210 29370
rect 2270 29310 2310 29370
rect 2370 29310 2410 29370
rect 2470 29310 2510 29370
rect 2570 29310 2610 29370
rect 2670 29310 2710 29370
rect 2770 29310 2810 29370
rect 2870 29310 2910 29370
rect 2970 29310 3010 29370
rect 3070 29310 3110 29370
rect 3170 29310 3210 29370
rect 3270 29310 3310 29370
rect 3370 29310 3410 29370
rect 3470 29310 3510 29370
rect 3570 29310 3610 29370
rect 3670 29310 3710 29370
rect 3770 29310 3810 29370
rect 3870 29310 3910 29370
rect 3970 29310 4010 29370
rect 4070 29310 4110 29370
rect 4170 29310 4210 29370
rect 4270 29310 4310 29370
rect 4370 29310 4410 29370
rect 4470 29310 4510 29370
rect 4570 29310 4610 29370
rect 4670 29310 4710 29370
rect 4770 29310 4810 29370
rect 4870 29310 4910 29370
rect 4970 29310 5010 29370
rect 5070 29310 5110 29370
rect 5170 29310 5210 29370
rect 5270 29310 5310 29370
rect 5370 29310 5410 29370
rect 5470 29310 5510 29370
rect 5570 29310 5610 29370
rect 5670 29310 5710 29370
rect 5770 29310 5810 29370
rect 5870 29310 5910 29370
rect 5970 29310 6010 29370
rect 6070 29310 6110 29370
rect 6170 29310 6210 29370
rect 6270 29310 6310 29370
rect 2170 29300 6310 29310
rect 7320 26610 20640 26620
rect 7320 26570 7360 26610
rect 7400 26570 7440 26610
rect 7480 26570 7520 26610
rect 7560 26570 7600 26610
rect 7640 26570 7680 26610
rect 7720 26570 7760 26610
rect 7800 26570 7840 26610
rect 7880 26570 7920 26610
rect 7960 26570 8000 26610
rect 8040 26570 8080 26610
rect 8120 26570 8160 26610
rect 8200 26570 8240 26610
rect 8280 26570 8320 26610
rect 8360 26570 8400 26610
rect 8440 26570 8480 26610
rect 8520 26570 8560 26610
rect 8600 26570 8640 26610
rect 8680 26570 8720 26610
rect 8760 26570 8800 26610
rect 8840 26570 8880 26610
rect 8920 26570 8960 26610
rect 9000 26570 9040 26610
rect 9080 26570 9120 26610
rect 9160 26570 9200 26610
rect 9240 26570 9280 26610
rect 9320 26570 9360 26610
rect 9400 26570 9440 26610
rect 9480 26570 9520 26610
rect 9560 26570 9600 26610
rect 9640 26570 9680 26610
rect 9720 26570 9760 26610
rect 9800 26570 9840 26610
rect 9880 26570 9920 26610
rect 9960 26570 10000 26610
rect 10040 26570 10080 26610
rect 10120 26570 10160 26610
rect 10200 26570 10240 26610
rect 10280 26570 10320 26610
rect 10360 26570 10400 26610
rect 10440 26570 10480 26610
rect 10520 26570 10560 26610
rect 10600 26570 10640 26610
rect 10680 26570 10720 26610
rect 10760 26570 10800 26610
rect 10840 26570 10880 26610
rect 10920 26570 10960 26610
rect 11000 26570 11040 26610
rect 11080 26570 11120 26610
rect 11160 26570 11200 26610
rect 11240 26570 11280 26610
rect 11320 26570 11360 26610
rect 11400 26570 11440 26610
rect 11480 26570 11520 26610
rect 11560 26570 11600 26610
rect 11640 26570 11680 26610
rect 11720 26570 11760 26610
rect 11800 26570 11840 26610
rect 11880 26570 11920 26610
rect 11960 26570 12000 26610
rect 12040 26570 12080 26610
rect 12120 26570 12160 26610
rect 12200 26570 12240 26610
rect 12280 26570 12320 26610
rect 12360 26570 12400 26610
rect 12440 26570 12480 26610
rect 12520 26570 12560 26610
rect 12600 26570 12640 26610
rect 12680 26570 12720 26610
rect 12760 26570 12800 26610
rect 12840 26570 12880 26610
rect 12920 26570 12960 26610
rect 13000 26570 13040 26610
rect 13080 26570 13120 26610
rect 13160 26570 13200 26610
rect 13240 26570 13280 26610
rect 13320 26570 13360 26610
rect 13400 26570 13440 26610
rect 13480 26570 13520 26610
rect 13560 26570 13600 26610
rect 13640 26570 13680 26610
rect 13720 26570 13760 26610
rect 13800 26570 13840 26610
rect 13880 26570 13920 26610
rect 13960 26570 14000 26610
rect 14040 26570 14080 26610
rect 14120 26570 14160 26610
rect 14200 26570 14240 26610
rect 14280 26570 14320 26610
rect 14360 26570 14400 26610
rect 14440 26570 14480 26610
rect 14520 26570 14560 26610
rect 14600 26570 14640 26610
rect 14680 26570 14720 26610
rect 14760 26570 14800 26610
rect 14840 26570 14880 26610
rect 14920 26570 14960 26610
rect 15000 26570 15040 26610
rect 15080 26570 15120 26610
rect 15160 26570 15200 26610
rect 15240 26570 15280 26610
rect 15320 26570 15360 26610
rect 15400 26570 15440 26610
rect 15480 26570 15520 26610
rect 15560 26570 15600 26610
rect 15640 26570 15680 26610
rect 15720 26570 15760 26610
rect 15800 26570 15840 26610
rect 15880 26570 15920 26610
rect 15960 26570 16000 26610
rect 16040 26570 16080 26610
rect 16120 26570 16160 26610
rect 16200 26570 16240 26610
rect 16280 26570 16320 26610
rect 16360 26570 16400 26610
rect 16440 26570 16480 26610
rect 16520 26570 16560 26610
rect 16600 26570 16640 26610
rect 16680 26570 16720 26610
rect 16760 26570 16800 26610
rect 16840 26570 16880 26610
rect 16920 26570 16960 26610
rect 17000 26570 17040 26610
rect 17080 26570 17120 26610
rect 17160 26570 17200 26610
rect 17240 26570 17280 26610
rect 17320 26570 17360 26610
rect 17400 26570 17440 26610
rect 17480 26570 17520 26610
rect 17560 26570 17600 26610
rect 17640 26570 17680 26610
rect 17720 26570 17760 26610
rect 17800 26570 17840 26610
rect 17880 26570 17920 26610
rect 17960 26570 18000 26610
rect 18040 26570 18080 26610
rect 18120 26570 18160 26610
rect 18200 26570 18240 26610
rect 18280 26570 18320 26610
rect 18360 26570 18400 26610
rect 18440 26570 18480 26610
rect 18520 26570 18560 26610
rect 18600 26570 18640 26610
rect 18680 26570 18720 26610
rect 18760 26570 18800 26610
rect 18840 26570 18880 26610
rect 18920 26570 18960 26610
rect 19000 26570 19040 26610
rect 19080 26570 19120 26610
rect 19160 26570 19200 26610
rect 19240 26570 19280 26610
rect 19320 26570 19360 26610
rect 19400 26570 19440 26610
rect 19480 26570 19520 26610
rect 19560 26570 19600 26610
rect 19640 26570 19680 26610
rect 19720 26570 19760 26610
rect 19800 26570 19840 26610
rect 19880 26570 19920 26610
rect 19960 26570 20000 26610
rect 20040 26570 20080 26610
rect 20120 26570 20160 26610
rect 20200 26570 20240 26610
rect 20280 26570 20320 26610
rect 20360 26570 20400 26610
rect 20440 26570 20480 26610
rect 20520 26570 20560 26610
rect 20600 26570 20640 26610
rect 7320 26560 20640 26570
rect 7280 21000 20640 21010
rect 7280 20960 7320 21000
rect 7360 20960 7400 21000
rect 7440 20960 7480 21000
rect 7520 20960 7560 21000
rect 7600 20960 7640 21000
rect 7680 20960 7720 21000
rect 7760 20960 7800 21000
rect 7840 20960 7880 21000
rect 7920 20960 7960 21000
rect 8000 20960 8040 21000
rect 8080 20960 8120 21000
rect 8160 20960 8200 21000
rect 8240 20960 8280 21000
rect 8320 20960 8360 21000
rect 8400 20960 8440 21000
rect 8480 20960 8520 21000
rect 8560 20960 8600 21000
rect 8640 20960 8680 21000
rect 8720 20960 8760 21000
rect 8800 20960 8840 21000
rect 8880 20960 8920 21000
rect 8960 20960 9000 21000
rect 9040 20960 9080 21000
rect 9120 20960 9160 21000
rect 9200 20960 9260 21000
rect 9300 20960 9340 21000
rect 9380 20960 9420 21000
rect 9460 20960 9500 21000
rect 9540 20960 9580 21000
rect 9620 20960 9660 21000
rect 9700 20960 9740 21000
rect 9780 20960 9820 21000
rect 9860 20960 9900 21000
rect 9940 20960 9980 21000
rect 10020 20960 10060 21000
rect 10100 20960 10140 21000
rect 10180 20960 10220 21000
rect 10260 20960 10300 21000
rect 10340 20960 10380 21000
rect 10420 20960 10460 21000
rect 10500 20960 10540 21000
rect 10580 20960 10620 21000
rect 10660 20960 10700 21000
rect 10740 20960 10780 21000
rect 10820 20960 10860 21000
rect 10900 20960 10940 21000
rect 10980 20960 11020 21000
rect 11060 20960 11100 21000
rect 11140 20960 11180 21000
rect 11220 20960 11260 21000
rect 11300 20960 11340 21000
rect 11380 20960 11420 21000
rect 11460 20960 11500 21000
rect 11540 20960 11580 21000
rect 11620 20960 11660 21000
rect 11700 20960 11740 21000
rect 11780 20960 11820 21000
rect 11860 20960 11900 21000
rect 11940 20960 11980 21000
rect 12020 20960 12060 21000
rect 12100 20960 12140 21000
rect 12180 20960 12220 21000
rect 12260 20960 12300 21000
rect 12340 20960 12380 21000
rect 12420 20960 12460 21000
rect 12500 20960 12540 21000
rect 12580 20960 12620 21000
rect 12660 20960 12700 21000
rect 12740 20960 12780 21000
rect 12820 20960 12880 21000
rect 12920 20960 12960 21000
rect 13000 20960 13040 21000
rect 13080 20960 13120 21000
rect 13160 20960 13200 21000
rect 13240 20960 13280 21000
rect 13320 20960 13360 21000
rect 13400 20960 13440 21000
rect 13480 20960 13520 21000
rect 13560 20960 13600 21000
rect 13640 20960 13680 21000
rect 13720 20960 13760 21000
rect 13800 20960 13840 21000
rect 13880 20960 13920 21000
rect 13960 20960 14000 21000
rect 14040 20960 14080 21000
rect 14120 20960 14160 21000
rect 14200 20960 14240 21000
rect 14280 20960 14320 21000
rect 14360 20960 14400 21000
rect 14440 20960 14480 21000
rect 14520 20960 14560 21000
rect 14600 20960 14640 21000
rect 14680 20960 14720 21000
rect 14760 20960 14800 21000
rect 14840 20960 14880 21000
rect 14920 20960 14960 21000
rect 15000 20960 15040 21000
rect 15080 20960 15120 21000
rect 15160 20960 15200 21000
rect 15240 20960 15280 21000
rect 15320 20960 15360 21000
rect 15400 20960 15440 21000
rect 15480 20960 15520 21000
rect 15560 20960 15600 21000
rect 15640 20960 15680 21000
rect 15720 20960 15760 21000
rect 15800 20960 15840 21000
rect 15880 20960 15920 21000
rect 15960 20960 16000 21000
rect 16040 20960 16080 21000
rect 16120 20960 16160 21000
rect 16200 20960 16240 21000
rect 16280 20960 16320 21000
rect 16360 20960 16400 21000
rect 16440 20960 16480 21000
rect 16520 20960 16560 21000
rect 16600 20960 16640 21000
rect 16680 20960 16720 21000
rect 16760 20960 16800 21000
rect 16840 20960 16880 21000
rect 16920 20960 16960 21000
rect 17000 20960 17040 21000
rect 17080 20960 17120 21000
rect 17160 20960 17200 21000
rect 17240 20960 17280 21000
rect 17320 20960 17360 21000
rect 17400 20960 17440 21000
rect 17480 20960 17520 21000
rect 17560 20960 17600 21000
rect 17640 20960 17680 21000
rect 17720 20960 17760 21000
rect 17800 20960 17840 21000
rect 17880 20960 17920 21000
rect 17960 20960 18000 21000
rect 18040 20960 18080 21000
rect 18120 20960 18160 21000
rect 18200 20960 18240 21000
rect 18280 20960 18320 21000
rect 18360 20960 18400 21000
rect 18440 20960 18480 21000
rect 18520 20960 18560 21000
rect 18600 20960 18640 21000
rect 18680 20960 18720 21000
rect 18760 20960 18800 21000
rect 18840 20960 18880 21000
rect 18920 20960 18960 21000
rect 19000 20960 19040 21000
rect 19080 20960 19120 21000
rect 19160 20960 19200 21000
rect 19240 20960 19280 21000
rect 19320 20960 19360 21000
rect 19400 20960 19440 21000
rect 19480 20960 19520 21000
rect 19560 20960 19600 21000
rect 19640 20960 19680 21000
rect 19720 20960 19760 21000
rect 19800 20960 19840 21000
rect 19880 20960 19920 21000
rect 19960 20960 20000 21000
rect 20040 20960 20080 21000
rect 20120 20960 20160 21000
rect 20200 20960 20240 21000
rect 20280 20960 20320 21000
rect 20360 20960 20400 21000
rect 20440 20960 20480 21000
rect 20520 20960 20560 21000
rect 20600 20960 20640 21000
rect 7280 20950 20640 20960
rect 7280 20470 8230 20480
rect 7280 20430 7320 20470
rect 7360 20430 7400 20470
rect 7440 20430 7480 20470
rect 7520 20430 7560 20470
rect 7600 20430 7640 20470
rect 7680 20430 7720 20470
rect 7760 20430 7800 20470
rect 7840 20430 7880 20470
rect 7920 20430 7960 20470
rect 8000 20430 8040 20470
rect 8080 20430 8120 20470
rect 8160 20430 8230 20470
rect 7280 20420 8230 20430
rect 8310 20020 20640 20030
rect 8310 19980 8360 20020
rect 8400 19980 8440 20020
rect 8480 19980 8520 20020
rect 8560 19980 8600 20020
rect 8640 19980 8680 20020
rect 8720 19980 8760 20020
rect 8800 19980 8840 20020
rect 8880 19980 8920 20020
rect 8960 19980 9000 20020
rect 9040 19980 9080 20020
rect 9120 19980 9160 20020
rect 9200 19980 9260 20020
rect 9300 19980 9340 20020
rect 9380 19980 9420 20020
rect 9460 19980 9500 20020
rect 9540 19980 9580 20020
rect 9620 19980 9660 20020
rect 9700 19980 9740 20020
rect 9780 19980 9820 20020
rect 9860 19980 9900 20020
rect 9940 19980 9980 20020
rect 10020 19980 10060 20020
rect 10100 19980 10140 20020
rect 10180 19980 10220 20020
rect 10260 19980 10300 20020
rect 10340 19980 10380 20020
rect 10420 19980 10460 20020
rect 10500 19980 10540 20020
rect 10580 19980 10620 20020
rect 10660 19980 10700 20020
rect 10740 19980 10780 20020
rect 10820 19980 10860 20020
rect 10900 19980 10940 20020
rect 10980 19980 11020 20020
rect 11060 19980 11100 20020
rect 11140 19980 11180 20020
rect 11220 19980 11260 20020
rect 11300 19980 11340 20020
rect 11380 19980 11420 20020
rect 11460 19980 11500 20020
rect 11540 19980 11580 20020
rect 11620 19980 11660 20020
rect 11700 19980 11740 20020
rect 11780 19980 11820 20020
rect 11860 19980 11900 20020
rect 11940 19980 11980 20020
rect 12020 19980 12060 20020
rect 12100 19980 12140 20020
rect 12180 19980 12220 20020
rect 12260 19980 12300 20020
rect 12340 19980 12380 20020
rect 12420 19980 12460 20020
rect 12500 19980 12540 20020
rect 12580 19980 12620 20020
rect 12660 19980 12700 20020
rect 12740 19980 12780 20020
rect 12820 19980 12860 20020
rect 12900 19980 12940 20020
rect 12980 19980 13040 20020
rect 13080 19980 13120 20020
rect 13160 19980 13200 20020
rect 13240 19980 13280 20020
rect 13320 19980 13360 20020
rect 13400 19980 13440 20020
rect 13480 19980 13520 20020
rect 13560 19980 13600 20020
rect 13640 19980 13680 20020
rect 13720 19980 13760 20020
rect 13800 19980 13840 20020
rect 13880 19980 13920 20020
rect 13960 19980 14000 20020
rect 14040 19980 14080 20020
rect 14120 19980 14160 20020
rect 14200 19980 14240 20020
rect 14280 19980 14320 20020
rect 14360 19980 14400 20020
rect 14440 19980 14480 20020
rect 14520 19980 14560 20020
rect 14600 19980 14640 20020
rect 14680 19980 14720 20020
rect 14760 19980 14800 20020
rect 14840 19980 14880 20020
rect 14920 19980 14960 20020
rect 15000 19980 15040 20020
rect 15080 19980 15120 20020
rect 15160 19980 15200 20020
rect 15240 19980 15280 20020
rect 15320 19980 15360 20020
rect 15400 19980 15440 20020
rect 15480 19980 15520 20020
rect 15560 19980 15600 20020
rect 15640 19980 15680 20020
rect 15720 19980 15760 20020
rect 15800 19980 15840 20020
rect 15880 19980 15920 20020
rect 15960 19980 16000 20020
rect 16040 19980 16080 20020
rect 16120 19980 16160 20020
rect 16200 19980 16240 20020
rect 16280 19980 16320 20020
rect 16360 19980 16400 20020
rect 16440 19980 16480 20020
rect 16520 19980 16560 20020
rect 16600 19980 16640 20020
rect 16680 19980 16720 20020
rect 16760 19980 16800 20020
rect 16840 19980 16880 20020
rect 16920 19980 16960 20020
rect 17000 19980 17040 20020
rect 17080 19980 17120 20020
rect 17160 19980 17200 20020
rect 17240 19980 17280 20020
rect 17320 19980 17360 20020
rect 17400 19980 17440 20020
rect 17480 19980 17520 20020
rect 17560 19980 17600 20020
rect 17640 19980 17680 20020
rect 17720 19980 17760 20020
rect 17800 19980 17840 20020
rect 17880 19980 17920 20020
rect 17960 19980 18000 20020
rect 18040 19980 18080 20020
rect 18120 19980 18160 20020
rect 18200 19980 18240 20020
rect 18280 19980 18320 20020
rect 18360 19980 18400 20020
rect 18440 19980 18480 20020
rect 18520 19980 18560 20020
rect 18600 19980 18640 20020
rect 18680 19980 18720 20020
rect 18760 19980 18800 20020
rect 18840 19980 18880 20020
rect 18920 19980 18960 20020
rect 19000 19980 19040 20020
rect 19080 19980 19120 20020
rect 19160 19980 19200 20020
rect 19240 19980 19280 20020
rect 19320 19980 19360 20020
rect 19400 19980 19440 20020
rect 19480 19980 19520 20020
rect 19560 19980 19600 20020
rect 19640 19980 19680 20020
rect 19720 19980 19760 20020
rect 19800 19980 19840 20020
rect 19880 19980 19920 20020
rect 19960 19980 20000 20020
rect 20040 19980 20080 20020
rect 20120 19980 20160 20020
rect 20200 19980 20240 20020
rect 20280 19980 20320 20020
rect 20360 19980 20400 20020
rect 20440 19980 20480 20020
rect 20520 19980 20560 20020
rect 20600 19980 20640 20020
rect 8310 19970 20640 19980
rect 9670 14340 21120 14350
rect 9670 14300 9700 14340
rect 9740 14300 9790 14340
rect 9830 14300 9870 14340
rect 9910 14300 9950 14340
rect 9990 14300 10030 14340
rect 10070 14300 10110 14340
rect 10150 14300 10190 14340
rect 10230 14300 10270 14340
rect 10310 14300 10350 14340
rect 10390 14300 10430 14340
rect 10470 14300 10510 14340
rect 10550 14300 10590 14340
rect 10630 14300 10670 14340
rect 10710 14300 10750 14340
rect 10790 14300 10830 14340
rect 10870 14300 10910 14340
rect 10950 14300 10990 14340
rect 11030 14300 11070 14340
rect 11110 14300 11150 14340
rect 11190 14300 11230 14340
rect 11270 14300 11310 14340
rect 11350 14300 11390 14340
rect 11430 14300 11470 14340
rect 11510 14300 11550 14340
rect 11590 14300 11630 14340
rect 11670 14300 11710 14340
rect 11750 14300 11790 14340
rect 11830 14300 11870 14340
rect 11910 14300 11950 14340
rect 11990 14300 12030 14340
rect 12070 14300 12110 14340
rect 12150 14300 12190 14340
rect 12230 14300 12270 14340
rect 12310 14300 12350 14340
rect 12390 14300 12430 14340
rect 12470 14300 12510 14340
rect 12550 14300 12590 14340
rect 12630 14300 12670 14340
rect 12710 14300 12750 14340
rect 12790 14300 12830 14340
rect 12870 14300 12910 14340
rect 12950 14300 12990 14340
rect 13030 14300 13070 14340
rect 13110 14300 13150 14340
rect 13230 14300 13270 14340
rect 13310 14300 13350 14340
rect 13390 14300 13430 14340
rect 13470 14300 13510 14340
rect 13550 14300 13590 14340
rect 13630 14300 13670 14340
rect 13710 14300 13750 14340
rect 13790 14300 13830 14340
rect 13870 14300 13910 14340
rect 13950 14300 13990 14340
rect 14030 14300 14070 14340
rect 14110 14300 14150 14340
rect 14190 14300 14230 14340
rect 14270 14300 14310 14340
rect 14350 14300 14390 14340
rect 14430 14300 14470 14340
rect 14510 14300 14550 14340
rect 14590 14300 14630 14340
rect 14670 14300 14710 14340
rect 14750 14300 14790 14340
rect 14830 14300 14870 14340
rect 14910 14300 14950 14340
rect 14990 14300 15030 14340
rect 15070 14300 15110 14340
rect 15150 14300 15190 14340
rect 15230 14300 15270 14340
rect 15310 14300 15350 14340
rect 15390 14300 15430 14340
rect 15470 14300 15510 14340
rect 15550 14300 15590 14340
rect 15630 14300 15670 14340
rect 15710 14300 15750 14340
rect 15790 14300 15830 14340
rect 15870 14300 15910 14340
rect 15950 14300 15990 14340
rect 16030 14300 16070 14340
rect 16110 14300 16150 14340
rect 16190 14300 16230 14340
rect 16270 14300 16310 14340
rect 16350 14300 16390 14340
rect 16430 14300 16470 14340
rect 16510 14300 16550 14340
rect 16590 14300 16630 14340
rect 16670 14300 16710 14340
rect 16750 14300 16790 14340
rect 16830 14300 16870 14340
rect 16910 14300 16950 14340
rect 16990 14300 17030 14340
rect 17070 14300 17110 14340
rect 17150 14300 17190 14340
rect 17230 14300 17270 14340
rect 17310 14300 17350 14340
rect 17390 14300 17430 14340
rect 17470 14300 17510 14340
rect 17550 14300 17590 14340
rect 17630 14300 17670 14340
rect 17710 14300 17750 14340
rect 17790 14300 17830 14340
rect 17870 14300 17910 14340
rect 17950 14300 17990 14340
rect 18030 14300 18070 14340
rect 18110 14300 18150 14340
rect 18190 14300 18230 14340
rect 18270 14300 18310 14340
rect 18350 14300 18390 14340
rect 18430 14300 18470 14340
rect 18510 14300 18550 14340
rect 18590 14300 18630 14340
rect 18670 14300 18710 14340
rect 18750 14300 18790 14340
rect 18830 14300 18870 14340
rect 18910 14300 18950 14340
rect 18990 14300 19030 14340
rect 19070 14300 19110 14340
rect 19150 14300 19190 14340
rect 19230 14300 19270 14340
rect 19310 14300 19350 14340
rect 19390 14300 19430 14340
rect 19470 14300 19510 14340
rect 19550 14300 19590 14340
rect 19630 14300 19670 14340
rect 19710 14300 19750 14340
rect 19790 14300 19830 14340
rect 19870 14300 19910 14340
rect 19950 14300 19990 14340
rect 20030 14300 20070 14340
rect 20110 14300 20150 14340
rect 20190 14300 20230 14340
rect 20270 14300 20310 14340
rect 20350 14300 20390 14340
rect 20430 14300 20470 14340
rect 20510 14300 20550 14340
rect 20590 14300 20630 14340
rect 20670 14300 20710 14340
rect 20750 14300 20790 14340
rect 20830 14300 20870 14340
rect 20910 14300 20950 14340
rect 20990 14300 21030 14340
rect 21070 14300 21120 14340
rect 9670 14290 21120 14300
rect 7280 13370 21110 13380
rect 7280 13330 7320 13370
rect 7360 13330 7400 13370
rect 7440 13330 7480 13370
rect 7520 13330 7560 13370
rect 7600 13330 7640 13370
rect 7680 13330 7720 13370
rect 7760 13330 7800 13370
rect 7840 13330 7880 13370
rect 7920 13330 7960 13370
rect 8000 13330 8040 13370
rect 8080 13330 8120 13370
rect 8160 13330 8200 13370
rect 8240 13330 8280 13370
rect 8320 13330 8360 13370
rect 8400 13330 8440 13370
rect 8480 13330 8520 13370
rect 8560 13330 8600 13370
rect 8640 13330 8680 13370
rect 8720 13330 8760 13370
rect 8800 13330 8840 13370
rect 8880 13330 8920 13370
rect 8960 13330 9000 13370
rect 9040 13330 9080 13370
rect 9120 13330 9160 13370
rect 9200 13330 9240 13370
rect 9280 13330 9320 13370
rect 9360 13330 9400 13370
rect 9440 13330 9480 13370
rect 9520 13330 9560 13370
rect 9600 13330 9640 13370
rect 9680 13330 9720 13370
rect 9760 13330 9800 13370
rect 9840 13330 9890 13370
rect 9930 13330 9970 13370
rect 10010 13330 10050 13370
rect 10090 13330 10130 13370
rect 10170 13330 10210 13370
rect 10250 13330 10290 13370
rect 10330 13330 10370 13370
rect 10410 13330 10450 13370
rect 10490 13330 10530 13370
rect 10570 13330 10610 13370
rect 10650 13330 10690 13370
rect 10730 13330 10770 13370
rect 10810 13330 10850 13370
rect 10890 13330 10930 13370
rect 10970 13330 11010 13370
rect 11050 13330 11090 13370
rect 11130 13330 11170 13370
rect 11210 13330 11250 13370
rect 11290 13330 11330 13370
rect 11370 13330 11410 13370
rect 11450 13330 11490 13370
rect 11530 13330 11570 13370
rect 11610 13330 11650 13370
rect 11690 13330 11730 13370
rect 11770 13330 11810 13370
rect 11850 13330 11890 13370
rect 11930 13330 11970 13370
rect 12010 13330 12050 13370
rect 12090 13330 12130 13370
rect 12170 13330 12210 13370
rect 12250 13330 12290 13370
rect 12330 13330 12370 13370
rect 12410 13330 12450 13370
rect 12490 13330 12530 13370
rect 12570 13330 12610 13370
rect 12650 13330 12690 13370
rect 12730 13330 12770 13370
rect 12810 13330 12850 13370
rect 12890 13330 12930 13370
rect 12970 13330 13010 13370
rect 13050 13330 13090 13370
rect 13130 13330 13170 13370
rect 13210 13330 13250 13370
rect 13290 13330 13330 13370
rect 13400 13330 13440 13370
rect 13480 13330 13520 13370
rect 13560 13330 13600 13370
rect 13640 13330 13680 13370
rect 13720 13330 13760 13370
rect 13800 13330 13840 13370
rect 13880 13330 13920 13370
rect 13960 13330 14000 13370
rect 14040 13330 14080 13370
rect 14120 13330 14160 13370
rect 14200 13330 14240 13370
rect 14280 13330 14320 13370
rect 14360 13330 14400 13370
rect 14440 13330 14480 13370
rect 14520 13330 14560 13370
rect 14600 13330 14640 13370
rect 14680 13330 14720 13370
rect 14760 13330 14800 13370
rect 14840 13330 14880 13370
rect 14920 13330 14960 13370
rect 15000 13330 15040 13370
rect 15080 13330 15120 13370
rect 15160 13330 15200 13370
rect 15240 13330 15280 13370
rect 15320 13330 15360 13370
rect 15400 13330 15440 13370
rect 15480 13330 15520 13370
rect 15560 13330 15600 13370
rect 15640 13330 15680 13370
rect 15720 13330 15760 13370
rect 15800 13330 15840 13370
rect 15880 13330 15920 13370
rect 15960 13330 16000 13370
rect 16040 13330 16080 13370
rect 16120 13330 16160 13370
rect 16200 13330 16240 13370
rect 16280 13330 16320 13370
rect 16360 13330 16400 13370
rect 16440 13330 16480 13370
rect 16520 13330 16560 13370
rect 16600 13330 16640 13370
rect 16680 13330 16720 13370
rect 16760 13330 16800 13370
rect 16840 13330 16880 13370
rect 16920 13330 16960 13370
rect 17000 13330 17040 13370
rect 17080 13330 17120 13370
rect 17160 13330 17200 13370
rect 17240 13330 17280 13370
rect 17320 13330 17360 13370
rect 17400 13330 17440 13370
rect 17480 13330 17520 13370
rect 17560 13330 17600 13370
rect 17640 13330 17680 13370
rect 17720 13330 17760 13370
rect 17800 13330 17840 13370
rect 17880 13330 17920 13370
rect 17960 13330 18000 13370
rect 18040 13330 18080 13370
rect 18120 13330 18160 13370
rect 18200 13330 18240 13370
rect 18280 13330 18320 13370
rect 18360 13330 18400 13370
rect 18440 13330 18480 13370
rect 18520 13330 18560 13370
rect 18600 13330 18640 13370
rect 18680 13330 18720 13370
rect 18760 13330 18800 13370
rect 18840 13330 18880 13370
rect 18920 13330 18960 13370
rect 19000 13330 19040 13370
rect 19080 13330 19120 13370
rect 19160 13330 19200 13370
rect 19240 13330 19280 13370
rect 19320 13330 19360 13370
rect 19400 13330 19440 13370
rect 19480 13330 19520 13370
rect 19560 13330 19600 13370
rect 19640 13330 19680 13370
rect 19720 13330 19760 13370
rect 19800 13330 19840 13370
rect 19880 13330 19920 13370
rect 19960 13330 20000 13370
rect 20040 13330 20080 13370
rect 20120 13330 20160 13370
rect 20200 13330 20240 13370
rect 20280 13330 20320 13370
rect 20360 13330 20400 13370
rect 20440 13330 20480 13370
rect 20520 13330 20560 13370
rect 20600 13330 20640 13370
rect 20680 13330 20720 13370
rect 20760 13330 20800 13370
rect 20840 13330 20880 13370
rect 20920 13330 20960 13370
rect 21000 13330 21040 13370
rect 21080 13330 21110 13370
rect 7280 13320 21110 13330
rect 7280 9720 7790 9730
rect 8470 9720 21120 9730
rect 7280 9680 7320 9720
rect 7360 9680 7400 9720
rect 7440 9680 7480 9720
rect 7520 9680 7560 9720
rect 7600 9680 7640 9720
rect 7680 9680 7720 9720
rect 7760 9680 7790 9720
rect 7280 9670 7790 9680
rect 7710 9650 7790 9670
rect 8470 9680 8520 9720
rect 8560 9680 8600 9720
rect 8640 9680 8680 9720
rect 8720 9680 8760 9720
rect 8800 9680 8840 9720
rect 8880 9680 8920 9720
rect 8960 9680 9000 9720
rect 9040 9680 9080 9720
rect 9120 9680 9160 9720
rect 9200 9680 9240 9720
rect 9280 9680 9320 9720
rect 9360 9680 9400 9720
rect 9440 9680 9480 9720
rect 9520 9680 9560 9720
rect 9600 9680 9640 9720
rect 9680 9680 9720 9720
rect 9760 9680 9800 9720
rect 9840 9680 9890 9720
rect 9930 9680 9970 9720
rect 10010 9680 10050 9720
rect 10090 9680 10130 9720
rect 10170 9680 10210 9720
rect 10250 9680 10290 9720
rect 10330 9680 10370 9720
rect 10410 9680 10450 9720
rect 10490 9680 10530 9720
rect 10570 9680 10610 9720
rect 10650 9680 10690 9720
rect 10730 9680 10770 9720
rect 10810 9680 10850 9720
rect 10890 9680 10930 9720
rect 10970 9680 11010 9720
rect 11050 9680 11090 9720
rect 11130 9680 11170 9720
rect 11210 9680 11250 9720
rect 11290 9680 11330 9720
rect 11370 9680 11410 9720
rect 11450 9680 11490 9720
rect 11530 9680 11570 9720
rect 11610 9680 11650 9720
rect 11690 9680 11730 9720
rect 11770 9680 11810 9720
rect 11850 9680 11890 9720
rect 11930 9680 11970 9720
rect 12010 9680 12050 9720
rect 12090 9680 12130 9720
rect 12170 9680 12210 9720
rect 12250 9680 12290 9720
rect 12330 9680 12370 9720
rect 12410 9680 12450 9720
rect 12490 9680 12530 9720
rect 12570 9680 12610 9720
rect 12650 9680 12690 9720
rect 12730 9680 12770 9720
rect 12810 9680 12850 9720
rect 12890 9680 12930 9720
rect 12970 9680 13010 9720
rect 13050 9680 13090 9720
rect 13130 9680 13170 9720
rect 13210 9680 13250 9720
rect 13290 9680 13330 9720
rect 13370 9680 13410 9720
rect 13450 9680 13490 9720
rect 13530 9680 13570 9720
rect 13610 9680 13650 9720
rect 13690 9680 13730 9720
rect 13770 9680 13810 9720
rect 13850 9680 13890 9720
rect 13930 9680 13970 9720
rect 14010 9680 14050 9720
rect 14090 9680 14130 9720
rect 14170 9680 14210 9720
rect 14250 9680 14290 9720
rect 14330 9680 14370 9720
rect 14410 9680 14450 9720
rect 14490 9680 14530 9720
rect 14570 9680 14610 9720
rect 14650 9680 14690 9720
rect 14730 9680 14770 9720
rect 14810 9680 14850 9720
rect 14890 9680 14930 9720
rect 14970 9680 15010 9720
rect 15050 9680 15090 9720
rect 15130 9680 15170 9720
rect 15210 9680 15250 9720
rect 15290 9680 15330 9720
rect 15370 9680 15410 9720
rect 15450 9680 15490 9720
rect 15530 9680 15570 9720
rect 15610 9680 15650 9720
rect 15690 9680 15730 9720
rect 15770 9680 15810 9720
rect 15850 9680 15890 9720
rect 15930 9680 15970 9720
rect 16010 9680 16050 9720
rect 16090 9680 16130 9720
rect 16170 9680 16210 9720
rect 16250 9680 16290 9720
rect 16330 9680 16370 9720
rect 16410 9680 16450 9720
rect 16490 9680 16530 9720
rect 16570 9680 16610 9720
rect 16650 9680 16690 9720
rect 16730 9680 16770 9720
rect 16810 9680 16850 9720
rect 16890 9680 16930 9720
rect 16970 9680 17010 9720
rect 17050 9680 17090 9720
rect 17130 9680 17170 9720
rect 17210 9680 17250 9720
rect 17290 9680 17330 9720
rect 17370 9680 17410 9720
rect 17450 9680 17490 9720
rect 17530 9680 17570 9720
rect 17610 9680 17650 9720
rect 17690 9680 17730 9720
rect 17770 9680 17810 9720
rect 17850 9680 17890 9720
rect 17930 9680 17970 9720
rect 18010 9680 18050 9720
rect 18090 9680 18130 9720
rect 18170 9680 18210 9720
rect 18250 9680 18290 9720
rect 18330 9680 18370 9720
rect 18410 9680 18450 9720
rect 18490 9680 18530 9720
rect 18570 9680 18610 9720
rect 18650 9680 18690 9720
rect 18730 9680 18770 9720
rect 18810 9680 18850 9720
rect 18890 9680 18930 9720
rect 18970 9680 19010 9720
rect 19050 9680 19090 9720
rect 19130 9680 19170 9720
rect 19210 9680 19250 9720
rect 19290 9680 19330 9720
rect 19370 9680 19410 9720
rect 19450 9680 19490 9720
rect 19530 9680 19570 9720
rect 19610 9680 19650 9720
rect 19690 9680 19730 9720
rect 19770 9680 19810 9720
rect 19850 9680 19890 9720
rect 19930 9680 19970 9720
rect 20010 9680 20050 9720
rect 20090 9680 20130 9720
rect 20170 9680 20210 9720
rect 20250 9680 20290 9720
rect 20330 9680 20370 9720
rect 20410 9680 20450 9720
rect 20490 9680 20530 9720
rect 20570 9680 20610 9720
rect 20650 9680 20690 9720
rect 20730 9680 20770 9720
rect 20810 9680 20850 9720
rect 20890 9680 20930 9720
rect 20970 9680 21010 9720
rect 21050 9680 21120 9720
rect 8470 9670 21120 9680
rect 8470 9650 8530 9670
rect 7710 9630 8530 9650
rect 7710 9590 7740 9630
rect 7780 9590 7820 9630
rect 7860 9590 7900 9630
rect 7940 9590 7980 9630
rect 8020 9590 8060 9630
rect 8100 9590 8140 9630
rect 8180 9590 8220 9630
rect 8260 9590 8300 9630
rect 8340 9590 8380 9630
rect 8420 9590 8460 9630
rect 8500 9590 8530 9630
rect 7710 9570 8530 9590
rect 12100 6990 12160 7000
rect 9870 6980 17060 6990
rect 9870 6930 9900 6980
rect 9960 6930 10120 6980
rect 10180 6930 10340 6980
rect 10400 6930 10560 6980
rect 10620 6930 10780 6980
rect 10840 6930 11000 6980
rect 11060 6930 11220 6980
rect 11280 6930 11440 6980
rect 11500 6930 11660 6980
rect 11720 6930 11880 6980
rect 11940 6930 12100 6980
rect 12160 6930 12320 6980
rect 12380 6930 12540 6980
rect 12600 6930 12760 6980
rect 12820 6930 12980 6980
rect 13040 6930 13200 6980
rect 13260 6930 13670 6980
rect 13730 6930 13890 6980
rect 13950 6930 14110 6980
rect 14170 6930 14330 6980
rect 14390 6930 14550 6980
rect 14610 6930 14770 6980
rect 14830 6930 14990 6980
rect 15050 6930 15210 6980
rect 15270 6930 15430 6980
rect 15490 6930 15650 6980
rect 15710 6930 15870 6980
rect 15930 6930 16090 6980
rect 16150 6930 16310 6980
rect 16370 6930 16530 6980
rect 16590 6930 16750 6980
rect 16810 6930 16970 6980
rect 17030 6930 17060 6980
rect 9870 6920 17060 6930
rect 13600 5990 17020 6000
rect 13600 5940 13630 5990
rect 13690 5940 13850 5990
rect 13910 5940 14070 5990
rect 14130 5940 14290 5990
rect 14350 5940 14510 5990
rect 14570 5940 14730 5990
rect 14790 5940 14950 5990
rect 15010 5940 15170 5990
rect 15230 5940 15390 5990
rect 15450 5940 15610 5990
rect 15670 5940 15830 5990
rect 15890 5940 16050 5990
rect 16110 5940 16270 5990
rect 16330 5940 16490 5990
rect 16550 5940 16710 5990
rect 16770 5940 16930 5990
rect 16990 5940 17020 5990
rect 13600 5930 17020 5940
rect 15830 5920 15890 5930
rect 9870 5870 13170 5880
rect 9870 5830 9930 5870
rect 9970 5830 10010 5870
rect 10050 5830 10090 5870
rect 10130 5830 10170 5870
rect 10210 5830 10250 5870
rect 10290 5830 10330 5870
rect 10370 5830 10410 5870
rect 10450 5830 10490 5870
rect 10530 5830 10610 5870
rect 10650 5830 10690 5870
rect 10730 5830 10770 5870
rect 10810 5830 10850 5870
rect 10890 5830 10930 5870
rect 10970 5830 11010 5870
rect 11050 5830 11090 5870
rect 11130 5830 11170 5870
rect 11210 5830 11250 5870
rect 11290 5830 11370 5870
rect 11410 5830 11450 5870
rect 11490 5830 11530 5870
rect 11570 5830 11610 5870
rect 11650 5830 11690 5870
rect 11730 5830 11770 5870
rect 11810 5830 11850 5870
rect 11890 5830 11930 5870
rect 11970 5830 12010 5870
rect 12050 5830 12130 5870
rect 12170 5830 12210 5870
rect 12250 5830 12290 5870
rect 12330 5830 12370 5870
rect 12410 5830 12450 5870
rect 12490 5830 12530 5870
rect 12570 5830 12610 5870
rect 12650 5830 12690 5870
rect 12730 5830 12770 5870
rect 12810 5830 12850 5870
rect 12890 5830 12930 5870
rect 12970 5830 13010 5870
rect 13050 5830 13090 5870
rect 13130 5830 13170 5870
rect 9870 5820 13170 5830
<< psubdiffcont >>
rect 3089 41640 3169 41680
rect 21620 41090 21680 41160
rect 21720 41090 21780 41160
rect 21830 41090 21890 41160
rect 21930 41090 21990 41160
rect 22030 41090 22090 41160
rect 22130 41090 22190 41160
rect 22230 41090 22290 41160
rect 22330 41090 22390 41160
rect 22430 41090 22490 41160
rect 22530 41090 22590 41160
rect 22630 41090 22690 41160
rect 22730 41090 22790 41160
rect 22830 41090 22890 41160
rect 22930 41090 22990 41160
rect 23030 41090 23090 41160
rect 23130 41090 23190 41160
rect 23230 41090 23290 41160
rect 23330 41090 23390 41160
rect 23430 41090 23490 41160
rect 23530 41090 23590 41160
rect 6009 40850 6070 40910
rect 2649 39500 2709 39560
rect 2749 39500 2809 39560
rect 2849 39500 2909 39560
rect 2949 39500 3009 39560
rect 3049 39500 3109 39560
rect 3149 39500 3209 39560
rect 3249 39500 3309 39560
rect 3349 39500 3409 39560
rect 3449 39500 3509 39560
rect 3549 39500 3609 39560
rect 3649 39500 3709 39560
rect 3749 39500 3809 39560
rect 3849 39500 3909 39560
rect 3949 39500 4009 39560
rect 4049 39500 4109 39560
rect 4149 39500 4209 39560
rect 4249 39500 4309 39560
rect 4349 39500 4409 39560
rect 4449 39500 4509 39560
rect 4549 39500 4609 39560
rect 4649 39500 4709 39560
rect 4749 39500 4809 39560
rect 4849 39500 4909 39560
rect 4949 39500 5009 39560
rect 5049 39500 5109 39560
rect 5149 39500 5209 39560
rect 5249 39500 5309 39560
rect 6349 39500 6409 39560
rect 6449 39500 6509 39560
rect 6549 39500 6609 39560
rect 6649 39500 6709 39560
rect 6749 39500 6809 39560
rect 6849 39500 6909 39560
rect 6949 39500 7009 39560
rect 7049 39500 7109 39560
rect 7149 39500 7209 39560
rect 7249 39500 7309 39560
rect 7349 39500 7409 39560
rect 7479 39500 7539 39560
rect 7579 39500 7639 39560
rect 7679 39500 7739 39560
rect 7779 39500 7839 39560
rect 7879 39500 7939 39560
rect 7979 39500 8039 39560
rect 8079 39500 8139 39560
rect 8179 39500 8239 39560
rect 8279 39500 8339 39560
rect 8379 39500 8439 39560
rect 8479 39500 8539 39560
rect 8629 39500 8689 39560
rect 8729 39500 8789 39560
rect 8829 39500 8889 39560
rect 8929 39500 8989 39560
rect 9029 39500 9089 39560
rect 9129 39500 9189 39560
rect 9229 39500 9289 39560
rect 9329 39500 9389 39560
rect 9429 39500 9489 39560
rect 9529 39500 9589 39560
rect 9629 39500 9689 39560
rect 9739 39500 9799 39560
rect 9839 39500 9899 39560
rect 3810 37120 3870 37180
rect 3910 37120 3970 37180
rect 4010 37120 4070 37180
rect 4110 37120 4170 37180
rect 4210 37120 4270 37180
rect 4310 37120 4370 37180
rect 4410 37120 4470 37180
rect 4510 37120 4570 37180
rect 4610 37120 4670 37180
rect 4710 37120 4770 37180
rect 4810 37120 4870 37180
rect 4910 37120 4970 37180
rect 5010 37120 5070 37180
rect 5110 37120 5170 37180
rect 5210 37120 5270 37180
rect 5310 37120 5370 37180
rect 5410 37120 5470 37180
rect 5510 37120 5570 37180
rect 5610 37120 5670 37180
rect 5710 37120 5770 37180
rect 5810 37120 5870 37180
rect 5910 37120 5970 37180
rect 6010 37120 6070 37180
rect 6110 37120 6170 37180
rect 6380 36660 6440 36720
rect 6480 36660 6540 36720
rect 6580 36660 6640 36720
rect 6680 36660 6740 36720
rect 6780 36660 6840 36720
rect 6880 36660 6940 36720
rect 6980 36660 7040 36720
rect 7080 36660 7140 36720
rect 7180 36660 7240 36720
rect 7280 36660 7340 36720
rect 7380 36660 7440 36720
rect 7480 36660 7540 36720
rect 7580 36660 7640 36720
rect 7680 36660 7740 36720
rect 7780 36660 7840 36720
rect 7880 36660 7940 36720
rect 7980 36660 8040 36720
rect 8080 36660 8140 36720
rect 8180 36660 8240 36720
rect 8280 36660 8340 36720
rect 8380 36660 8440 36720
rect 8480 36660 8540 36720
rect 8580 36660 8640 36720
rect 8680 36660 8740 36720
rect 8780 36660 8840 36720
rect 8880 36660 8940 36720
rect 8980 36660 9040 36720
rect 9080 36660 9140 36720
rect 9180 36660 9240 36720
rect 9280 36660 9340 36720
rect 9380 36660 9440 36720
rect 9480 36660 9540 36720
rect 9580 36660 9640 36720
rect 9680 36660 9740 36720
rect 9780 36660 9840 36720
rect 9880 36660 9940 36720
rect 9980 36660 10040 36720
rect 10080 36660 10140 36720
rect 10180 36660 10240 36720
rect 10280 36660 10340 36720
rect 10380 36660 10440 36720
rect 10480 36660 10540 36720
rect 10580 36660 10640 36720
rect 10680 36660 10740 36720
rect 10780 36660 10840 36720
rect 15790 35570 15900 35630
rect 16510 34130 16570 34200
rect 16610 34130 16670 34200
rect 16710 34130 16770 34200
rect 16810 34130 16870 34200
rect 16910 34130 16970 34200
rect 17010 34130 17070 34200
rect 17110 34130 17170 34200
rect 17210 34130 17270 34200
rect 17310 34130 17370 34200
rect 17410 34130 17470 34200
rect 17510 34130 17570 34200
rect 17610 34130 17670 34200
rect 17710 34130 17770 34200
rect 17810 34130 17870 34200
rect 17910 34130 17970 34200
rect 18010 34130 18070 34200
rect 18110 34130 18170 34200
rect 18210 34130 18270 34200
rect 18310 34130 18370 34200
rect 18410 34130 18470 34200
rect 18510 34130 18570 34200
rect 18610 34130 18670 34200
rect 18710 34130 18770 34200
rect 18810 34130 18870 34200
rect 18910 34130 18970 34200
rect 19010 34130 19070 34200
rect 19110 34130 19170 34200
rect 19210 34130 19270 34200
rect 19310 34130 19370 34200
rect 19410 34130 19470 34200
rect 19510 34130 19570 34200
rect 19610 34130 19670 34200
rect 19710 34130 19770 34200
rect 19810 34130 19870 34200
rect 19910 34130 19970 34200
rect 20010 34130 20070 34200
rect 20110 34130 20170 34200
rect 20210 34130 20270 34200
rect 20310 34130 20370 34200
rect 20410 34130 20470 34200
rect 20510 34130 20570 34200
rect 20610 34130 20670 34200
rect 20710 34130 20770 34200
rect 20810 34130 20870 34200
rect 20910 34130 20970 34200
rect 21010 34130 21070 34200
rect 21110 34130 21170 34200
rect 21210 34130 21270 34200
rect 21310 34130 21370 34200
rect 21410 34130 21470 34200
rect 21510 34130 21570 34200
rect 21610 34130 21670 34200
rect 21710 34130 21770 34200
rect 21810 34130 21870 34200
rect 21910 34130 21970 34200
rect 22010 34130 22070 34200
rect 22110 34130 22170 34200
rect 22210 34130 22270 34200
rect 22310 34130 22370 34200
rect 22410 34130 22470 34200
rect 22510 34130 22570 34200
rect 22610 34130 22670 34200
rect 22710 34130 22770 34200
rect 22810 34130 22870 34200
rect 22910 34130 22970 34200
rect 23010 34130 23070 34200
rect 23110 34130 23170 34200
rect 23210 34130 23270 34200
rect 23310 34130 23370 34200
rect 23410 34130 23470 34200
rect 23510 34130 23570 34200
rect 23620 34130 23680 34200
rect 23720 34130 23780 34200
rect 23820 34130 23880 34200
rect 23920 34130 23980 34200
rect 24020 34130 24080 34200
rect 24120 34130 24180 34200
rect 24220 34130 24280 34200
rect 24320 34130 24380 34200
rect 24420 34130 24480 34200
rect 24520 34130 24580 34200
rect 24620 34130 24680 34200
rect 24720 34130 24780 34200
rect 24820 34130 24880 34200
rect 24920 34130 24980 34200
rect 25020 34130 25080 34200
rect 25120 34130 25180 34200
rect 25220 34130 25280 34200
rect 25320 34130 25380 34200
rect 14400 31950 14510 32010
rect 2210 31670 2270 31730
rect 2310 31670 2370 31730
rect 2410 31670 2470 31730
rect 2510 31670 2570 31730
rect 2610 31670 2670 31730
rect 2710 31670 2770 31730
rect 2810 31670 2870 31730
rect 2910 31670 2970 31730
rect 3010 31670 3070 31730
rect 3110 31670 3170 31730
rect 3210 31670 3270 31730
rect 3310 31670 3370 31730
rect 3410 31670 3470 31730
rect 3510 31670 3570 31730
rect 3610 31670 3670 31730
rect 3710 31670 3770 31730
rect 3810 31670 3870 31730
rect 3910 31670 3970 31730
rect 4010 31670 4070 31730
rect 4110 31670 4170 31730
rect 4210 31670 4270 31730
rect 4310 31670 4370 31730
rect 4410 31670 4470 31730
rect 4510 31670 4570 31730
rect 4610 31670 4670 31730
rect 4710 31670 4770 31730
rect 4810 31670 4870 31730
rect 4910 31670 4970 31730
rect 5010 31670 5070 31730
rect 5110 31670 5170 31730
rect 5210 31670 5270 31730
rect 5310 31670 5370 31730
rect 5410 31670 5470 31730
rect 5510 31670 5570 31730
rect 5610 31670 5670 31730
rect 5710 31670 5770 31730
rect 5810 31670 5870 31730
rect 5910 31670 5970 31730
rect 6010 31670 6070 31730
rect 6110 31670 6170 31730
rect 6210 31670 6270 31730
rect 6470 31320 6530 31380
rect 6580 31320 6640 31380
rect 6690 31320 6750 31380
rect 6800 31320 6860 31380
rect 6910 31320 6970 31380
rect 7020 31320 7080 31380
rect 7130 31320 7190 31380
rect 7240 31320 7300 31380
rect 7350 31320 7410 31380
rect 7460 31320 7520 31380
rect 7570 31320 7630 31380
rect 7680 31320 7740 31380
rect 7790 31320 7850 31380
rect 7900 31320 7960 31380
rect 8010 31320 8070 31380
rect 8120 31320 8180 31380
rect 8230 31320 8290 31380
rect 8340 31320 8400 31380
rect 8450 31320 8510 31380
rect 8560 31320 8620 31380
rect 8670 31320 8730 31380
rect 8780 31320 8840 31380
rect 8890 31320 8950 31380
rect 9000 31320 9060 31380
rect 9110 31320 9170 31380
rect 9220 31320 9280 31380
rect 9330 31320 9390 31380
rect 9440 31320 9500 31380
rect 9550 31320 9610 31380
rect 9660 31320 9720 31380
rect 9770 31320 9830 31380
rect 9880 31320 9940 31380
rect 9990 31320 10050 31380
rect 10100 31320 10160 31380
rect 10210 31320 10270 31380
rect 10320 31320 10380 31380
rect 10430 31320 10490 31380
rect 10540 31320 10600 31380
rect 10650 31320 10710 31380
rect 10760 31320 10820 31380
rect 10880 31320 10940 31380
rect 10990 31320 11050 31380
rect 11100 31320 11160 31380
rect 14870 30060 14930 30130
rect 14970 30060 15030 30130
rect 15070 30060 15130 30130
rect 15170 30060 15230 30130
rect 15270 30060 15330 30130
rect 15370 30060 15430 30130
rect 15470 30060 15530 30130
rect 15570 30060 15630 30130
rect 15670 30060 15730 30130
rect 15780 30060 15840 30130
rect 15880 30060 15940 30130
rect 15990 30060 16050 30130
rect 16130 30060 16190 30130
rect 16270 30060 16330 30130
rect 16370 30060 16430 30130
rect 16470 30060 16530 30130
rect 16570 30060 16630 30130
rect 16670 30060 16730 30130
rect 16770 30060 16830 30130
rect 16870 30060 16930 30130
rect 16970 30060 17030 30130
rect 17070 30060 17130 30130
rect 17170 30060 17230 30130
rect 17270 30060 17330 30130
rect 17370 30060 17430 30130
rect 17470 30060 17530 30130
rect 17570 30060 17630 30130
rect 17670 30060 17730 30130
rect 17770 30060 17830 30130
rect 17870 30060 17930 30130
rect 17970 30060 18030 30130
rect 18070 30060 18130 30130
rect 18170 30060 18230 30130
rect 18270 30060 18330 30130
rect 18370 30060 18430 30130
rect 18470 30060 18530 30130
rect 18570 30060 18630 30130
rect 18670 30060 18730 30130
rect 18770 30060 18830 30130
rect 18870 30060 18930 30130
rect 18970 30060 19030 30130
rect 19070 30060 19130 30130
rect 19170 30060 19230 30130
rect 19270 30060 19330 30130
rect 19370 30060 19430 30130
rect 19470 30060 19530 30130
rect 19570 30060 19630 30130
rect 19670 30060 19730 30130
rect 19770 30060 19830 30130
rect 19870 30060 19930 30130
rect 19970 30060 20030 30130
rect 20070 30060 20130 30130
rect 20170 30060 20230 30130
rect 20270 30060 20330 30130
rect 20370 30060 20430 30130
rect 20470 30060 20530 30130
rect 20570 30060 20630 30130
rect 20670 30060 20730 30130
rect 20770 30060 20830 30130
rect 20870 30060 20930 30130
rect 20970 30060 21030 30130
rect 21070 30060 21130 30130
rect 21170 30060 21230 30130
rect 21270 30060 21330 30130
rect 21370 30060 21430 30130
rect 21470 30060 21530 30130
rect 21570 30060 21630 30130
rect 21670 30060 21730 30130
rect 21770 30060 21830 30130
rect 21870 30060 21930 30130
rect 21970 30060 22030 30130
rect 22070 30060 22130 30130
rect 22170 30060 22230 30130
rect 22270 30060 22330 30130
rect 22370 30060 22430 30130
rect 22470 30060 22530 30130
rect 22570 30060 22630 30130
rect 22670 30060 22730 30130
rect 22770 30060 22830 30130
rect 22870 30060 22930 30130
rect 22970 30060 23030 30130
rect 23070 30060 23130 30130
rect 23170 30060 23230 30130
rect 23270 30060 23330 30130
rect 23370 30060 23430 30130
rect 23470 30060 23530 30130
rect 23570 30060 23630 30130
rect 23670 30060 23730 30130
rect 23770 30060 23830 30130
rect 23870 30060 23930 30130
rect 23970 30060 24030 30130
rect 24070 30060 24130 30130
rect 24170 30060 24230 30130
rect 24270 30060 24330 30130
rect 24370 30060 24430 30130
rect 24470 30060 24530 30130
rect 24570 30060 24630 30130
rect 24670 30060 24730 30130
rect 24770 30060 24830 30130
rect 24870 30060 24930 30130
rect 24970 30060 25030 30130
rect 25070 30060 25130 30130
rect 25170 30060 25230 30130
rect 25270 30060 25330 30130
rect 25370 30060 25430 30130
rect 25470 30060 25530 30130
rect 25570 30060 25630 30130
rect 7320 24250 7360 24290
rect 7400 24250 7440 24290
rect 7480 24250 7520 24290
rect 7560 24250 7600 24290
rect 7640 24250 7680 24290
rect 7720 24250 7760 24290
rect 7800 24250 7840 24290
rect 7890 24250 7930 24290
rect 7970 24250 8010 24290
rect 8050 24250 8090 24290
rect 8130 24250 8170 24290
rect 8210 24250 8250 24290
rect 8290 24250 8330 24290
rect 8400 24250 8440 24290
rect 8520 24250 8560 24290
rect 8600 24250 8640 24290
rect 8680 24250 8720 24290
rect 8760 24250 8800 24290
rect 8840 24250 8880 24290
rect 8920 24250 8960 24290
rect 9000 24250 9040 24290
rect 9080 24250 9120 24290
rect 9160 24250 9200 24290
rect 9270 24250 9310 24290
rect 9350 24250 9390 24290
rect 9430 24250 9470 24290
rect 9510 24250 9550 24290
rect 9590 24250 9630 24290
rect 9670 24250 9710 24290
rect 9750 24250 9790 24290
rect 9830 24250 9870 24290
rect 9910 24250 9950 24290
rect 9990 24250 10030 24290
rect 10070 24250 10110 24290
rect 10150 24250 10190 24290
rect 10230 24250 10270 24290
rect 10310 24250 10350 24290
rect 10390 24250 10430 24290
rect 10470 24250 10510 24290
rect 10550 24250 10590 24290
rect 10630 24250 10670 24290
rect 10710 24250 10750 24290
rect 10790 24250 10830 24290
rect 10870 24250 10910 24290
rect 10950 24250 10990 24290
rect 11030 24250 11070 24290
rect 11110 24250 11150 24290
rect 11190 24250 11230 24290
rect 11270 24250 11310 24290
rect 11350 24250 11390 24290
rect 11430 24250 11470 24290
rect 11510 24250 11550 24290
rect 11590 24250 11630 24290
rect 11670 24250 11710 24290
rect 11750 24250 11790 24290
rect 11830 24250 11870 24290
rect 11910 24250 11950 24290
rect 11990 24250 12030 24290
rect 12070 24250 12110 24290
rect 12150 24250 12190 24290
rect 12230 24250 12270 24290
rect 12310 24250 12350 24290
rect 12390 24250 12430 24290
rect 12470 24250 12510 24290
rect 12550 24250 12590 24290
rect 12630 24250 12670 24290
rect 12710 24250 12750 24290
rect 12790 24250 12830 24290
rect 12870 24250 12910 24290
rect 12950 24250 12990 24290
rect 13030 24250 13070 24290
rect 13110 24250 13150 24290
rect 13190 24250 13230 24290
rect 13270 24250 13310 24290
rect 13350 24250 13390 24290
rect 13430 24250 13470 24290
rect 13510 24250 13550 24290
rect 13590 24250 13630 24290
rect 13670 24250 13710 24290
rect 13750 24250 13790 24290
rect 13830 24250 13870 24290
rect 13910 24250 13950 24290
rect 13990 24250 14030 24290
rect 14070 24250 14110 24290
rect 14150 24250 14190 24290
rect 14230 24250 14270 24290
rect 14310 24250 14350 24290
rect 14390 24250 14430 24290
rect 14470 24250 14510 24290
rect 14550 24250 14590 24290
rect 14630 24250 14670 24290
rect 14710 24250 14750 24290
rect 14790 24250 14830 24290
rect 14870 24250 14910 24290
rect 14950 24250 14990 24290
rect 15030 24250 15070 24290
rect 15110 24250 15150 24290
rect 15190 24250 15230 24290
rect 15270 24250 15310 24290
rect 15350 24250 15390 24290
rect 15430 24250 15470 24290
rect 15510 24250 15550 24290
rect 15590 24250 15630 24290
rect 15670 24250 15710 24290
rect 15750 24250 15790 24290
rect 15830 24250 15870 24290
rect 15910 24250 15950 24290
rect 15990 24250 16030 24290
rect 16070 24250 16110 24290
rect 16150 24250 16190 24290
rect 16230 24250 16270 24290
rect 16310 24250 16350 24290
rect 16390 24250 16430 24290
rect 16470 24250 16510 24290
rect 16550 24250 16590 24290
rect 16630 24250 16670 24290
rect 16710 24250 16750 24290
rect 16790 24250 16830 24290
rect 16870 24250 16910 24290
rect 16950 24250 16990 24290
rect 17030 24250 17070 24290
rect 17110 24250 17150 24290
rect 17190 24250 17230 24290
rect 17270 24250 17310 24290
rect 17350 24250 17390 24290
rect 17430 24250 17470 24290
rect 17510 24250 17550 24290
rect 17590 24250 17630 24290
rect 17670 24250 17710 24290
rect 17750 24250 17790 24290
rect 17830 24250 17870 24290
rect 17910 24250 17950 24290
rect 17990 24250 18030 24290
rect 18070 24250 18110 24290
rect 18150 24250 18190 24290
rect 18230 24250 18270 24290
rect 18310 24250 18350 24290
rect 18390 24250 18430 24290
rect 18470 24250 18510 24290
rect 18550 24250 18590 24290
rect 18630 24250 18670 24290
rect 18710 24250 18750 24290
rect 18790 24250 18830 24290
rect 18870 24250 18910 24290
rect 18950 24250 18990 24290
rect 19030 24250 19070 24290
rect 19110 24250 19150 24290
rect 19190 24250 19230 24290
rect 19270 24250 19310 24290
rect 19350 24250 19390 24290
rect 19430 24250 19470 24290
rect 19510 24250 19550 24290
rect 19590 24250 19630 24290
rect 19670 24250 19710 24290
rect 19750 24250 19790 24290
rect 19830 24250 19870 24290
rect 19910 24250 19950 24290
rect 19990 24250 20030 24290
rect 20070 24250 20110 24290
rect 20150 24250 20190 24290
rect 20230 24250 20270 24290
rect 20310 24250 20350 24290
rect 20390 24250 20430 24290
rect 20470 24250 20510 24290
rect 20550 24250 20590 24290
rect 7310 23280 7350 23320
rect 7390 23280 7430 23320
rect 7470 23280 7510 23320
rect 7550 23280 7590 23320
rect 7630 23280 7670 23320
rect 7710 23280 7750 23320
rect 7790 23280 7830 23320
rect 7870 23280 7910 23320
rect 7950 23280 7990 23320
rect 8030 23280 8070 23320
rect 8110 23280 8150 23320
rect 8190 23280 8230 23320
rect 8270 23280 8310 23320
rect 8350 23280 8390 23320
rect 8430 23280 8470 23320
rect 8520 23280 8560 23320
rect 8600 23280 8640 23320
rect 8680 23280 8720 23320
rect 8760 23280 8800 23320
rect 8840 23280 8880 23320
rect 8920 23280 8960 23320
rect 9000 23280 9040 23320
rect 9080 23280 9120 23320
rect 9160 23280 9200 23320
rect 9270 23280 9310 23320
rect 9350 23280 9390 23320
rect 9430 23280 9470 23320
rect 9510 23280 9550 23320
rect 9590 23280 9630 23320
rect 9670 23280 9710 23320
rect 9750 23280 9790 23320
rect 9830 23280 9870 23320
rect 9910 23280 9950 23320
rect 9990 23280 10030 23320
rect 10070 23280 10110 23320
rect 10150 23280 10190 23320
rect 10230 23280 10270 23320
rect 10310 23280 10350 23320
rect 10390 23280 10430 23320
rect 10470 23280 10510 23320
rect 10550 23280 10590 23320
rect 10630 23280 10670 23320
rect 10710 23280 10750 23320
rect 10790 23280 10830 23320
rect 10870 23280 10910 23320
rect 10950 23280 10990 23320
rect 11030 23280 11070 23320
rect 11110 23280 11150 23320
rect 11190 23280 11230 23320
rect 11270 23280 11310 23320
rect 11350 23280 11390 23320
rect 11430 23280 11470 23320
rect 11510 23280 11550 23320
rect 11590 23280 11630 23320
rect 11670 23280 11710 23320
rect 11750 23280 11790 23320
rect 11830 23280 11870 23320
rect 11910 23280 11950 23320
rect 11990 23280 12030 23320
rect 12070 23280 12110 23320
rect 12150 23280 12190 23320
rect 12230 23280 12270 23320
rect 12310 23280 12350 23320
rect 12390 23280 12430 23320
rect 12470 23280 12510 23320
rect 12550 23280 12590 23320
rect 12630 23280 12670 23320
rect 12710 23280 12750 23320
rect 12790 23280 12830 23320
rect 12870 23280 12910 23320
rect 12950 23280 12990 23320
rect 13030 23280 13070 23320
rect 13110 23280 13150 23320
rect 13190 23280 13230 23320
rect 13270 23280 13310 23320
rect 13350 23280 13390 23320
rect 13430 23280 13470 23320
rect 13510 23280 13550 23320
rect 13590 23280 13630 23320
rect 13670 23280 13710 23320
rect 13750 23280 13790 23320
rect 13830 23280 13870 23320
rect 13910 23280 13950 23320
rect 13990 23280 14030 23320
rect 14070 23280 14110 23320
rect 14150 23280 14190 23320
rect 14230 23280 14270 23320
rect 14310 23280 14350 23320
rect 14390 23280 14430 23320
rect 14470 23280 14510 23320
rect 14550 23280 14590 23320
rect 14630 23280 14670 23320
rect 14710 23280 14750 23320
rect 14790 23280 14830 23320
rect 14870 23280 14910 23320
rect 14950 23280 14990 23320
rect 15030 23280 15070 23320
rect 15110 23280 15150 23320
rect 15190 23280 15230 23320
rect 15270 23280 15310 23320
rect 15350 23280 15390 23320
rect 15430 23280 15470 23320
rect 15510 23280 15550 23320
rect 15590 23280 15630 23320
rect 15670 23280 15710 23320
rect 15750 23280 15790 23320
rect 15830 23280 15870 23320
rect 15910 23280 15950 23320
rect 15990 23280 16030 23320
rect 16070 23280 16110 23320
rect 16150 23280 16190 23320
rect 16230 23280 16270 23320
rect 16310 23280 16350 23320
rect 16390 23280 16430 23320
rect 16470 23280 16510 23320
rect 16550 23280 16590 23320
rect 16630 23280 16670 23320
rect 16710 23280 16750 23320
rect 16790 23280 16830 23320
rect 16870 23280 16910 23320
rect 16950 23280 16990 23320
rect 17030 23280 17070 23320
rect 17110 23280 17150 23320
rect 17190 23280 17230 23320
rect 17270 23280 17310 23320
rect 17350 23280 17390 23320
rect 17430 23280 17470 23320
rect 17510 23280 17550 23320
rect 17590 23280 17630 23320
rect 17670 23280 17710 23320
rect 17750 23280 17790 23320
rect 17830 23280 17870 23320
rect 17910 23280 17950 23320
rect 17990 23280 18030 23320
rect 18070 23280 18110 23320
rect 18150 23280 18190 23320
rect 18230 23280 18270 23320
rect 18310 23280 18350 23320
rect 18390 23280 18430 23320
rect 18470 23280 18510 23320
rect 18550 23280 18590 23320
rect 18630 23280 18670 23320
rect 18710 23280 18750 23320
rect 18790 23280 18830 23320
rect 18870 23280 18910 23320
rect 18950 23280 18990 23320
rect 19030 23280 19070 23320
rect 19110 23280 19150 23320
rect 19190 23280 19230 23320
rect 19270 23280 19310 23320
rect 19350 23280 19390 23320
rect 19430 23280 19470 23320
rect 19510 23280 19550 23320
rect 19590 23280 19630 23320
rect 19670 23280 19710 23320
rect 19750 23280 19790 23320
rect 19830 23280 19870 23320
rect 19910 23280 19950 23320
rect 19990 23280 20030 23320
rect 20070 23280 20110 23320
rect 20150 23280 20190 23320
rect 20230 23280 20270 23320
rect 20310 23280 20350 23320
rect 20390 23280 20430 23320
rect 20470 23280 20510 23320
rect 20550 23280 20590 23320
rect 7320 17660 7360 17700
rect 7400 17660 7440 17700
rect 7480 17660 7520 17700
rect 7560 17660 7600 17700
rect 7640 17660 7680 17700
rect 7720 17660 7760 17700
rect 7800 17660 7840 17700
rect 7880 17660 7920 17700
rect 7960 17660 8000 17700
rect 8040 17660 8080 17700
rect 8120 17660 8160 17700
rect 8200 17660 8240 17700
rect 8280 17660 8320 17700
rect 8360 17660 8400 17700
rect 8440 17660 8480 17700
rect 8520 17660 8560 17700
rect 8600 17660 8640 17700
rect 8680 17660 8720 17700
rect 8760 17660 8800 17700
rect 8840 17660 8880 17700
rect 8920 17660 8960 17700
rect 9000 17660 9040 17700
rect 9080 17660 9120 17700
rect 9160 17660 9200 17700
rect 9270 17660 9310 17700
rect 9350 17660 9390 17700
rect 9430 17660 9470 17700
rect 9510 17660 9550 17700
rect 9590 17660 9630 17700
rect 9670 17660 9710 17700
rect 9750 17660 9790 17700
rect 9830 17660 9870 17700
rect 9910 17660 9950 17700
rect 9990 17660 10030 17700
rect 10070 17660 10110 17700
rect 10150 17660 10190 17700
rect 10230 17660 10270 17700
rect 10310 17660 10350 17700
rect 10390 17660 10430 17700
rect 10470 17660 10510 17700
rect 10550 17660 10590 17700
rect 10630 17660 10670 17700
rect 10710 17660 10750 17700
rect 10790 17660 10830 17700
rect 10870 17660 10910 17700
rect 10950 17660 10990 17700
rect 11030 17660 11070 17700
rect 11110 17660 11150 17700
rect 11190 17660 11230 17700
rect 11270 17660 11310 17700
rect 11350 17660 11390 17700
rect 11430 17660 11470 17700
rect 11510 17660 11550 17700
rect 11590 17660 11630 17700
rect 11670 17660 11710 17700
rect 11750 17660 11790 17700
rect 11830 17660 11870 17700
rect 11910 17660 11950 17700
rect 11990 17660 12030 17700
rect 12070 17660 12110 17700
rect 12150 17660 12190 17700
rect 12230 17660 12270 17700
rect 12310 17660 12350 17700
rect 12390 17660 12430 17700
rect 12470 17660 12510 17700
rect 12550 17660 12590 17700
rect 12630 17660 12670 17700
rect 12710 17660 12750 17700
rect 12790 17660 12830 17700
rect 12870 17660 12910 17700
rect 12950 17660 12990 17700
rect 13030 17660 13070 17700
rect 13110 17660 13150 17700
rect 13190 17660 13230 17700
rect 13270 17660 13310 17700
rect 13350 17660 13390 17700
rect 13430 17660 13470 17700
rect 13510 17660 13550 17700
rect 13590 17660 13630 17700
rect 13670 17660 13710 17700
rect 13750 17660 13790 17700
rect 13830 17660 13870 17700
rect 13910 17660 13950 17700
rect 13990 17660 14030 17700
rect 14070 17660 14110 17700
rect 14150 17660 14190 17700
rect 14230 17660 14270 17700
rect 14310 17660 14350 17700
rect 14390 17660 14430 17700
rect 14470 17660 14510 17700
rect 14550 17660 14590 17700
rect 14630 17660 14670 17700
rect 14710 17660 14750 17700
rect 14790 17660 14830 17700
rect 14870 17660 14910 17700
rect 14950 17660 14990 17700
rect 15030 17660 15070 17700
rect 15110 17660 15150 17700
rect 15190 17660 15230 17700
rect 15270 17660 15310 17700
rect 15350 17660 15390 17700
rect 15430 17660 15470 17700
rect 15510 17660 15550 17700
rect 15590 17660 15630 17700
rect 15670 17660 15710 17700
rect 15750 17660 15790 17700
rect 15830 17660 15870 17700
rect 15910 17660 15950 17700
rect 15990 17660 16030 17700
rect 16070 17660 16110 17700
rect 16150 17660 16190 17700
rect 16230 17660 16270 17700
rect 16310 17660 16350 17700
rect 16390 17660 16430 17700
rect 16470 17660 16510 17700
rect 16550 17660 16590 17700
rect 16630 17660 16670 17700
rect 16710 17660 16750 17700
rect 16790 17660 16830 17700
rect 16870 17660 16910 17700
rect 16950 17660 16990 17700
rect 17030 17660 17070 17700
rect 17110 17660 17150 17700
rect 17190 17660 17230 17700
rect 17270 17660 17310 17700
rect 17350 17660 17390 17700
rect 17430 17660 17470 17700
rect 17510 17660 17550 17700
rect 17590 17660 17630 17700
rect 17670 17660 17710 17700
rect 17750 17660 17790 17700
rect 17830 17660 17870 17700
rect 17910 17660 17950 17700
rect 17990 17660 18030 17700
rect 18070 17660 18110 17700
rect 18150 17660 18190 17700
rect 18230 17660 18270 17700
rect 18310 17660 18350 17700
rect 18390 17660 18430 17700
rect 18470 17660 18510 17700
rect 18550 17660 18590 17700
rect 18630 17660 18670 17700
rect 18710 17660 18750 17700
rect 18790 17660 18830 17700
rect 18870 17660 18910 17700
rect 18950 17660 18990 17700
rect 19030 17660 19070 17700
rect 19110 17660 19150 17700
rect 19190 17660 19230 17700
rect 19270 17660 19310 17700
rect 19350 17660 19390 17700
rect 19430 17660 19470 17700
rect 19510 17660 19550 17700
rect 19590 17660 19630 17700
rect 19670 17660 19710 17700
rect 19750 17660 19790 17700
rect 19830 17660 19870 17700
rect 19910 17660 19950 17700
rect 19990 17660 20030 17700
rect 20070 17660 20110 17700
rect 20150 17660 20190 17700
rect 20230 17660 20270 17700
rect 20310 17660 20350 17700
rect 20390 17660 20430 17700
rect 20470 17660 20510 17700
rect 20550 17660 20590 17700
rect 9710 15620 9750 15660
rect 9790 15620 9830 15660
rect 9870 15620 9910 15660
rect 9950 15620 9990 15660
rect 10030 15620 10070 15660
rect 10110 15620 10150 15660
rect 10190 15620 10230 15660
rect 10270 15620 10310 15660
rect 10350 15620 10390 15660
rect 10430 15620 10470 15660
rect 10510 15620 10550 15660
rect 10590 15620 10630 15660
rect 10670 15620 10710 15660
rect 10750 15620 10790 15660
rect 10830 15620 10870 15660
rect 10910 15620 10950 15660
rect 10990 15620 11030 15660
rect 11070 15620 11110 15660
rect 11150 15620 11190 15660
rect 11230 15620 11270 15660
rect 11310 15620 11350 15660
rect 11390 15620 11430 15660
rect 11470 15620 11510 15660
rect 11550 15620 11590 15660
rect 11630 15620 11670 15660
rect 11710 15620 11750 15660
rect 11790 15620 11830 15660
rect 11870 15620 11910 15660
rect 11950 15620 11990 15660
rect 12030 15620 12070 15660
rect 12110 15620 12150 15660
rect 12190 15620 12230 15660
rect 12270 15620 12310 15660
rect 12350 15620 12390 15660
rect 12430 15620 12470 15660
rect 12510 15620 12550 15660
rect 12590 15620 12630 15660
rect 12670 15620 12710 15660
rect 12750 15620 12790 15660
rect 12830 15620 12870 15660
rect 12910 15620 12950 15660
rect 12990 15620 13030 15660
rect 13070 15620 13110 15660
rect 13150 15620 13190 15660
rect 13230 15620 13270 15660
rect 13310 15620 13350 15660
rect 13390 15620 13430 15660
rect 13470 15620 13510 15660
rect 13550 15620 13590 15660
rect 13630 15620 13670 15660
rect 13710 15620 13750 15660
rect 13790 15620 13830 15660
rect 13870 15620 13910 15660
rect 13950 15620 13990 15660
rect 14030 15620 14070 15660
rect 14110 15620 14150 15660
rect 14190 15620 14230 15660
rect 14270 15620 14310 15660
rect 14350 15620 14390 15660
rect 14430 15620 14470 15660
rect 14510 15620 14550 15660
rect 14590 15620 14630 15660
rect 14670 15620 14710 15660
rect 14750 15620 14790 15660
rect 14830 15620 14870 15660
rect 14910 15620 14950 15660
rect 14990 15620 15030 15660
rect 15070 15620 15110 15660
rect 15150 15620 15190 15660
rect 15230 15620 15270 15660
rect 15310 15620 15350 15660
rect 15390 15620 15430 15660
rect 15470 15620 15510 15660
rect 15550 15620 15590 15660
rect 15630 15620 15670 15660
rect 15710 15620 15750 15660
rect 15790 15620 15830 15660
rect 15870 15620 15910 15660
rect 15950 15620 15990 15660
rect 16030 15620 16070 15660
rect 16110 15620 16150 15660
rect 16190 15620 16230 15660
rect 16270 15620 16310 15660
rect 16350 15620 16390 15660
rect 16430 15620 16470 15660
rect 16510 15620 16550 15660
rect 16590 15620 16630 15660
rect 16670 15620 16710 15660
rect 16750 15620 16790 15660
rect 16830 15620 16870 15660
rect 16910 15620 16950 15660
rect 16990 15620 17030 15660
rect 17070 15620 17110 15660
rect 17150 15620 17190 15660
rect 17230 15620 17270 15660
rect 17310 15620 17350 15660
rect 17390 15620 17430 15660
rect 17470 15620 17510 15660
rect 17550 15620 17590 15660
rect 17630 15620 17670 15660
rect 17710 15620 17750 15660
rect 17790 15620 17830 15660
rect 17870 15620 17910 15660
rect 17950 15620 17990 15660
rect 18030 15620 18070 15660
rect 18110 15620 18150 15660
rect 18190 15620 18230 15660
rect 18270 15620 18310 15660
rect 18350 15620 18390 15660
rect 18430 15620 18470 15660
rect 18510 15620 18550 15660
rect 18590 15620 18630 15660
rect 18670 15620 18710 15660
rect 18750 15620 18790 15660
rect 18830 15620 18870 15660
rect 18910 15620 18950 15660
rect 18990 15620 19030 15660
rect 19070 15620 19110 15660
rect 19150 15620 19190 15660
rect 19230 15620 19270 15660
rect 19310 15620 19350 15660
rect 19390 15620 19430 15660
rect 19470 15620 19510 15660
rect 19550 15620 19590 15660
rect 19630 15620 19670 15660
rect 19710 15620 19750 15660
rect 19800 15620 19840 15660
rect 19880 15620 19920 15660
rect 19960 15620 20000 15660
rect 20040 15620 20080 15660
rect 20120 15620 20160 15660
rect 20200 15620 20240 15660
rect 20280 15620 20320 15660
rect 20370 15620 20410 15660
rect 20450 15620 20490 15660
rect 20530 15620 20570 15660
rect 20610 15620 20650 15660
rect 20690 15620 20730 15660
rect 20770 15620 20810 15660
rect 20850 15620 20890 15660
rect 20930 15620 20970 15660
rect 21010 15620 21050 15660
rect 21090 15620 21130 15660
rect 9810 12010 9850 12050
rect 9890 12010 9930 12050
rect 9970 12010 10010 12050
rect 10050 12010 10090 12050
rect 10130 12010 10170 12050
rect 10210 12010 10250 12050
rect 10290 12010 10330 12050
rect 10370 12010 10410 12050
rect 10450 12010 10490 12050
rect 10530 12010 10570 12050
rect 10610 12010 10650 12050
rect 10690 12010 10730 12050
rect 10770 12010 10810 12050
rect 10850 12010 10890 12050
rect 10930 12010 10970 12050
rect 11010 12010 11050 12050
rect 11090 12010 11130 12050
rect 11170 12010 11210 12050
rect 11250 12010 11290 12050
rect 11330 12010 11370 12050
rect 11410 12010 11450 12050
rect 11490 12010 11530 12050
rect 11570 12010 11610 12050
rect 11650 12010 11690 12050
rect 11730 12010 11770 12050
rect 11810 12010 11850 12050
rect 11890 12010 11930 12050
rect 11970 12010 12010 12050
rect 12050 12010 12090 12050
rect 12130 12010 12170 12050
rect 12210 12010 12250 12050
rect 12290 12010 12330 12050
rect 12370 12010 12410 12050
rect 12450 12010 12490 12050
rect 12530 12010 12570 12050
rect 12610 12010 12650 12050
rect 12690 12010 12730 12050
rect 12770 12010 12810 12050
rect 12850 12010 12890 12050
rect 12930 12010 12970 12050
rect 13010 12010 13050 12050
rect 13090 12010 13130 12050
rect 13170 12010 13210 12050
rect 13250 12010 13290 12050
rect 13330 12010 13440 12050
rect 13480 12010 13520 12050
rect 13560 12010 13600 12050
rect 13640 12010 13680 12050
rect 13720 12010 13760 12050
rect 13800 12010 13840 12050
rect 13880 12010 13920 12050
rect 13960 12010 14000 12050
rect 14040 12010 14080 12050
rect 14120 12010 14160 12050
rect 14200 12010 14240 12050
rect 14280 12010 14320 12050
rect 14360 12010 14400 12050
rect 14440 12010 14480 12050
rect 14520 12010 14560 12050
rect 14600 12010 14640 12050
rect 14680 12010 14720 12050
rect 14760 12010 14800 12050
rect 14840 12010 14880 12050
rect 14920 12010 14960 12050
rect 15000 12010 15040 12050
rect 15080 12010 15120 12050
rect 15160 12010 15200 12050
rect 15240 12010 15280 12050
rect 15320 12010 15360 12050
rect 15400 12010 15440 12050
rect 15480 12010 15520 12050
rect 15560 12010 15600 12050
rect 15640 12010 15680 12050
rect 15720 12010 15760 12050
rect 15800 12010 15840 12050
rect 15880 12010 15920 12050
rect 15960 12010 16000 12050
rect 16040 12010 16080 12050
rect 16120 12010 16160 12050
rect 16200 12010 16240 12050
rect 16280 12010 16320 12050
rect 16360 12010 16400 12050
rect 16440 12010 16480 12050
rect 16520 12010 16560 12050
rect 16600 12010 16640 12050
rect 16680 12010 16720 12050
rect 16760 12010 16800 12050
rect 16840 12010 16880 12050
rect 16920 12010 16960 12050
rect 17000 12010 17040 12050
rect 17080 12010 17120 12050
rect 17160 12010 17200 12050
rect 17240 12010 17280 12050
rect 17320 12010 17360 12050
rect 17400 12010 17440 12050
rect 17480 12010 17520 12050
rect 17560 12010 17600 12050
rect 17640 12010 17680 12050
rect 17720 12010 17760 12050
rect 17800 12010 17840 12050
rect 17880 12010 17920 12050
rect 17960 12010 18000 12050
rect 18040 12010 18080 12050
rect 18120 12010 18160 12050
rect 18200 12010 18240 12050
rect 18280 12010 18320 12050
rect 18360 12010 18400 12050
rect 18440 12010 18480 12050
rect 18520 12010 18560 12050
rect 18600 12010 18640 12050
rect 18680 12010 18720 12050
rect 18760 12010 18800 12050
rect 18840 12010 18880 12050
rect 18920 12010 18960 12050
rect 19000 12010 19040 12050
rect 19080 12010 19120 12050
rect 19160 12010 19200 12050
rect 19240 12010 19280 12050
rect 19320 12010 19360 12050
rect 19400 12010 19440 12050
rect 19480 12010 19520 12050
rect 19560 12010 19600 12050
rect 19640 12010 19680 12050
rect 19720 12010 19760 12050
rect 19800 12010 19840 12050
rect 19890 12010 19930 12050
rect 19970 12010 20010 12050
rect 20050 12010 20090 12050
rect 20130 12010 20170 12050
rect 20210 12010 20250 12050
rect 20290 12010 20330 12050
rect 20370 12010 20410 12050
rect 20460 12010 20500 12050
rect 20540 12010 20580 12050
rect 20620 12010 20660 12050
rect 20700 12010 20740 12050
rect 20780 12010 20820 12050
rect 20860 12010 20900 12050
rect 20940 12010 20980 12050
rect 21020 12010 21060 12050
rect 7330 11960 7370 12000
rect 7410 11960 7450 12000
rect 7490 11960 7530 12000
rect 7570 11960 7610 12000
rect 7650 11960 7690 12000
rect 7730 11960 7770 12000
rect 7810 11960 7850 12000
rect 7890 11960 7930 12000
rect 7970 11960 8010 12000
rect 8050 11960 8090 12000
rect 8130 11960 8170 12000
rect 8210 11960 8250 12000
rect 8290 11960 8330 12000
rect 8370 11960 8410 12000
rect 8450 11960 8490 12000
rect 8530 11960 8570 12000
rect 8610 11960 8650 12000
rect 8690 11960 8730 12000
rect 8770 11960 8810 12000
rect 8850 11960 8890 12000
rect 8930 11960 8970 12000
rect 9010 11960 9050 12000
rect 9090 11960 9130 12000
rect 9170 11960 9210 12000
rect 9250 11960 9290 12000
rect 9330 11960 9370 12000
rect 9410 11960 9450 12000
rect 9490 11960 9530 12000
rect 9570 11960 9610 12000
rect 9650 11960 9690 12000
rect 9730 11960 9770 12000
rect 7720 11370 7760 11410
rect 7800 11370 7840 11410
rect 7880 11370 7920 11410
rect 7960 11370 8000 11410
rect 8040 11370 8080 11410
rect 8120 11370 8160 11410
rect 8200 11370 8240 11410
rect 8280 11370 8320 11410
rect 8360 11370 8400 11410
rect 8440 11370 8480 11410
rect 8520 11370 8560 11410
rect 7670 11290 7710 11330
rect 7670 11210 7710 11250
rect 7670 11130 7710 11170
rect 8550 11290 8590 11330
rect 8550 11210 8590 11250
rect 8550 11130 8590 11170
rect 7330 11050 7370 11090
rect 7410 11050 7450 11090
rect 7490 11050 7530 11090
rect 7570 11050 7610 11090
rect 7650 11050 7690 11090
rect 8610 11050 8650 11090
rect 8690 11050 8730 11090
rect 8770 11050 8810 11090
rect 8850 11050 8890 11090
rect 8930 11050 8970 11090
rect 9010 11050 9050 11090
rect 9090 11050 9130 11090
rect 9170 11050 9210 11090
rect 9250 11050 9290 11090
rect 9330 11050 9370 11090
rect 9410 11050 9450 11090
rect 9490 11050 9530 11090
rect 9570 11050 9610 11090
rect 9650 11050 9690 11090
rect 9730 11050 9770 11090
rect 9810 11000 9850 11040
rect 9890 11000 9930 11040
rect 9970 11000 10010 11040
rect 10050 11000 10090 11040
rect 10130 11000 10170 11040
rect 10210 11000 10250 11040
rect 10290 11000 10330 11040
rect 10370 11000 10410 11040
rect 10450 11000 10490 11040
rect 10530 11000 10570 11040
rect 10610 11000 10650 11040
rect 10690 11000 10730 11040
rect 10770 11000 10810 11040
rect 10850 11000 10890 11040
rect 10930 11000 10970 11040
rect 11010 11000 11050 11040
rect 11090 11000 11130 11040
rect 11170 11000 11210 11040
rect 11250 11000 11290 11040
rect 11330 11000 11370 11040
rect 11410 11000 11450 11040
rect 11490 11000 11530 11040
rect 11570 11000 11610 11040
rect 11650 11000 11690 11040
rect 11730 11000 11770 11040
rect 11810 11000 11850 11040
rect 11890 11000 11930 11040
rect 11970 11000 12010 11040
rect 12050 11000 12090 11040
rect 12130 11000 12170 11040
rect 12210 11000 12250 11040
rect 12290 11000 12330 11040
rect 12370 11000 12410 11040
rect 12450 11000 12490 11040
rect 12530 11000 12570 11040
rect 12610 11000 12650 11040
rect 12690 11000 12730 11040
rect 12770 11000 12810 11040
rect 12850 11000 12890 11040
rect 12930 11000 12970 11040
rect 13010 11000 13050 11040
rect 13090 11000 13130 11040
rect 13170 11000 13210 11040
rect 13250 11000 13290 11040
rect 13330 11000 13410 11040
rect 13450 11000 13490 11040
rect 13530 11000 13570 11040
rect 13610 11000 13650 11040
rect 13690 11000 13730 11040
rect 13770 11000 13810 11040
rect 13850 11000 13890 11040
rect 13930 11000 13970 11040
rect 14010 11000 14050 11040
rect 14090 11000 14130 11040
rect 14170 11000 14210 11040
rect 14250 11000 14290 11040
rect 14330 11000 14370 11040
rect 14410 11000 14450 11040
rect 14490 11000 14530 11040
rect 14570 11000 14610 11040
rect 14650 11000 14690 11040
rect 14730 11000 14770 11040
rect 14810 11000 14850 11040
rect 14890 11000 14930 11040
rect 14970 11000 15010 11040
rect 15050 11000 15090 11040
rect 15130 11000 15170 11040
rect 15210 11000 15250 11040
rect 15290 11000 15330 11040
rect 15370 11000 15410 11040
rect 15450 11000 15490 11040
rect 15530 11000 15570 11040
rect 15610 11000 15650 11040
rect 15690 11000 15730 11040
rect 15770 11000 15810 11040
rect 15850 11000 15890 11040
rect 15930 11000 15970 11040
rect 16010 11000 16050 11040
rect 16090 11000 16130 11040
rect 16170 11000 16210 11040
rect 16250 11000 16290 11040
rect 16330 11000 16370 11040
rect 16410 11000 16450 11040
rect 16490 11000 16530 11040
rect 16570 11000 16610 11040
rect 16650 11000 16690 11040
rect 16730 11000 16770 11040
rect 16810 11000 16850 11040
rect 16890 11000 16930 11040
rect 16970 11000 17010 11040
rect 17050 11000 17090 11040
rect 17130 11000 17170 11040
rect 17210 11000 17250 11040
rect 17290 11000 17330 11040
rect 17370 11000 17410 11040
rect 17450 11000 17490 11040
rect 17530 11000 17570 11040
rect 17610 11000 17650 11040
rect 17690 11000 17730 11040
rect 17770 11000 17810 11040
rect 17850 11000 17890 11040
rect 17930 11000 17970 11040
rect 18010 11000 18050 11040
rect 18090 11000 18130 11040
rect 18170 11000 18210 11040
rect 18250 11000 18290 11040
rect 18330 11000 18370 11040
rect 18410 11000 18450 11040
rect 18490 11000 18530 11040
rect 18570 11000 18610 11040
rect 18650 11000 18690 11040
rect 18730 11000 18770 11040
rect 18810 11000 18850 11040
rect 18890 11000 18930 11040
rect 18970 11000 19010 11040
rect 19050 11000 19090 11040
rect 19130 11000 19170 11040
rect 19210 11000 19250 11040
rect 19290 11000 19330 11040
rect 19370 11000 19410 11040
rect 19450 11000 19490 11040
rect 19540 11000 19580 11040
rect 19620 11000 19660 11040
rect 19700 11000 19740 11040
rect 19780 11000 19820 11040
rect 19860 11000 19900 11040
rect 19940 11000 19980 11040
rect 20020 11000 20060 11040
rect 20110 11000 20150 11040
rect 20190 11000 20230 11040
rect 20270 11000 20310 11040
rect 20350 11000 20390 11040
rect 20430 11000 20470 11040
rect 20510 11000 20550 11040
rect 20590 11000 20630 11040
rect 20670 11000 20710 11040
rect 20750 11000 20790 11040
rect 20830 11000 20870 11040
rect 20910 11000 20950 11040
rect 20990 11000 21030 11040
rect 21070 11000 21110 11040
rect 13630 2950 13690 3000
rect 13850 2950 13910 3000
rect 14070 2950 14130 3000
rect 14290 2950 14350 3000
rect 14510 2950 14570 3000
rect 14730 2950 14790 3000
rect 14950 2950 15010 3000
rect 15170 2950 15230 3000
rect 15390 2950 15450 3000
rect 15610 2950 15670 3000
rect 15830 2950 15890 3000
rect 16050 2950 16110 3000
rect 16270 2950 16330 3000
rect 16490 2950 16550 3000
rect 16710 2950 16770 3000
rect 24220 2660 24280 2720
rect 24220 2560 24280 2620
rect 24220 2460 24280 2520
rect 24220 2360 24280 2420
rect 24220 2260 24280 2320
rect 24220 2160 24280 2220
rect 24220 2060 24280 2120
rect 9890 1870 9950 1920
rect 10110 1870 10170 1920
rect 10330 1870 10390 1920
rect 10550 1870 10610 1920
rect 10770 1870 10830 1920
rect 10990 1870 11050 1920
rect 11210 1870 11270 1920
rect 11430 1870 11490 1920
rect 11650 1870 11710 1920
rect 11870 1870 11930 1920
rect 12090 1870 12150 1920
rect 12310 1870 12370 1920
rect 12530 1870 12590 1920
rect 12750 1870 12810 1920
rect 12970 1870 13030 1920
rect 13630 1870 13690 1920
rect 13850 1870 13910 1920
rect 14070 1870 14130 1920
rect 14290 1870 14350 1920
rect 14510 1870 14570 1920
rect 14730 1870 14790 1920
rect 14950 1870 15010 1920
rect 15170 1870 15230 1920
rect 15390 1870 15450 1920
rect 15610 1870 15670 1920
rect 15830 1870 15890 1920
rect 16050 1870 16110 1920
rect 16270 1870 16330 1920
rect 16490 1870 16550 1920
rect 16710 1870 16770 1920
<< nsubdiffcont >>
rect 21830 43280 21890 43350
rect 21930 43280 21990 43350
rect 22030 43280 22090 43350
rect 22130 43280 22190 43350
rect 22230 43280 22290 43350
rect 22330 43280 22390 43350
rect 22430 43280 22490 43350
rect 22530 43280 22590 43350
rect 22630 43280 22690 43350
rect 22730 43280 22790 43350
rect 22830 43280 22890 43350
rect 22930 43280 22990 43350
rect 23030 43280 23090 43350
rect 23130 43280 23190 43350
rect 23230 43280 23290 43350
rect 23330 43280 23390 43350
rect 23430 43280 23490 43350
rect 23530 43280 23590 43350
rect 2469 42110 2519 42160
rect 2559 42110 2609 42160
rect 2649 42110 2699 42160
rect 2739 42110 2789 42160
rect 2829 42110 2879 42160
rect 2919 42110 2969 42160
rect 3429 41900 3479 41950
rect 3519 41900 3569 41950
rect 3609 41900 3659 41950
rect 3699 41900 3749 41950
rect 3789 41900 3839 41950
rect 3879 41900 3929 41950
rect 3969 41900 4019 41950
rect 4059 41900 4109 41950
rect 4149 41900 4199 41950
rect 4239 41900 4289 41950
rect 4579 41890 4639 41950
rect 6009 41910 6069 41970
rect 6119 41910 6179 41970
rect 6229 41910 6289 41970
rect 6339 41910 6399 41970
rect 6449 41910 6509 41970
rect 6559 41910 6619 41970
rect 6669 41910 6729 41970
rect 6779 41910 6839 41970
rect 6889 41910 6949 41970
rect 6999 41910 7059 41970
rect 7109 41910 7169 41970
rect 7219 41910 7279 41970
rect 7329 41910 7389 41970
rect 7439 41910 7499 41970
rect 7549 41910 7609 41970
rect 7659 41910 7719 41970
rect 7769 41910 7829 41970
rect 7879 41910 7939 41970
rect 7989 41910 8049 41970
rect 8099 41910 8159 41970
rect 8209 41910 8269 41970
rect 8319 41910 8379 41970
rect 8429 41910 8489 41970
rect 8539 41910 8599 41970
rect 8649 41910 8709 41970
rect 8759 41910 8819 41970
rect 8869 41910 8929 41970
rect 8979 41910 9039 41970
rect 9089 41910 9149 41970
rect 9199 41910 9259 41970
rect 9309 41910 9369 41970
rect 9419 41910 9479 41970
rect 9529 41910 9589 41970
rect 9639 41910 9699 41970
rect 9749 41910 9809 41970
rect 9859 41910 9919 41970
rect 3320 40610 3380 40670
rect 3430 40610 3490 40670
rect 3540 40610 3600 40670
rect 3650 40610 3710 40670
rect 3760 40610 3820 40670
rect 3870 40610 3930 40670
rect 3980 40610 4040 40670
rect 4090 40610 4150 40670
rect 4659 40620 5399 40660
rect 6409 40590 6469 40650
rect 6519 40590 6579 40650
rect 6629 40590 6689 40650
rect 6739 40590 6799 40650
rect 6849 40590 6909 40650
rect 6959 40590 7019 40650
rect 7069 40590 7129 40650
rect 7179 40590 7239 40650
rect 7289 40590 7349 40650
rect 7399 40590 7459 40650
rect 7509 40590 7569 40650
rect 7619 40590 7679 40650
rect 7729 40590 7789 40650
rect 7839 40590 7899 40650
rect 7949 40590 8009 40650
rect 8059 40590 8119 40650
rect 8169 40590 8229 40650
rect 8279 40590 8339 40650
rect 8389 40590 8449 40650
rect 8499 40590 8559 40650
rect 8609 40590 8669 40650
rect 8719 40590 8779 40650
rect 8829 40590 8889 40650
rect 8939 40590 8999 40650
rect 9049 40590 9109 40650
rect 9159 40590 9219 40650
rect 9269 40590 9329 40650
rect 9379 40590 9439 40650
rect 9489 40590 9549 40650
rect 9599 40590 9659 40650
rect 9709 40590 9769 40650
rect 9819 40590 9879 40650
rect 15220 36270 15280 36340
rect 15320 36270 15380 36340
rect 15420 36270 15480 36340
rect 15520 36270 15580 36340
rect 15620 36270 15680 36340
rect 15720 36270 15780 36340
rect 15820 36270 15880 36340
rect 15920 36270 15980 36340
rect 16020 36270 16080 36340
rect 16120 36270 16180 36340
rect 16220 36270 16280 36340
rect 16320 36270 16380 36340
rect 16420 36270 16480 36340
rect 16520 36270 16580 36340
rect 16620 36270 16680 36340
rect 16720 36270 16780 36340
rect 16820 36270 16880 36340
rect 16920 36270 16980 36340
rect 17020 36270 17080 36340
rect 17120 36270 17180 36340
rect 17220 36270 17280 36340
rect 17320 36270 17380 36340
rect 17420 36270 17480 36340
rect 17520 36270 17580 36340
rect 17620 36270 17680 36340
rect 17720 36270 17780 36340
rect 17820 36270 17880 36340
rect 17920 36270 17980 36340
rect 18020 36270 18080 36340
rect 18120 36270 18180 36340
rect 18220 36270 18280 36340
rect 18320 36270 18380 36340
rect 18420 36270 18480 36340
rect 18520 36270 18580 36340
rect 18620 36270 18680 36340
rect 18720 36270 18780 36340
rect 18820 36270 18880 36340
rect 18920 36270 18980 36340
rect 19020 36270 19080 36340
rect 19120 36270 19180 36340
rect 19220 36270 19280 36340
rect 19320 36270 19380 36340
rect 19420 36270 19480 36340
rect 19520 36270 19580 36340
rect 19620 36270 19680 36340
rect 19720 36270 19780 36340
rect 19820 36270 19880 36340
rect 19920 36270 19980 36340
rect 20020 36270 20080 36340
rect 20120 36270 20180 36340
rect 20220 36270 20280 36340
rect 20320 36270 20380 36340
rect 20420 36270 20480 36340
rect 20520 36270 20580 36340
rect 20620 36270 20680 36340
rect 20720 36270 20780 36340
rect 20820 36270 20880 36340
rect 20920 36270 20980 36340
rect 21020 36270 21080 36340
rect 21120 36270 21180 36340
rect 21220 36270 21280 36340
rect 21320 36270 21380 36340
rect 21420 36270 21480 36340
rect 21520 36270 21580 36340
rect 21620 36270 21680 36340
rect 21720 36270 21780 36340
rect 21820 36270 21880 36340
rect 21920 36270 21980 36340
rect 22020 36270 22080 36340
rect 22120 36270 22180 36340
rect 22220 36270 22280 36340
rect 22320 36270 22380 36340
rect 22420 36270 22480 36340
rect 22520 36270 22580 36340
rect 22620 36270 22680 36340
rect 22720 36270 22780 36340
rect 22820 36270 22880 36340
rect 22920 36270 22980 36340
rect 23020 36270 23080 36340
rect 23120 36270 23180 36340
rect 23220 36270 23280 36340
rect 23320 36270 23380 36340
rect 23420 36270 23480 36340
rect 23520 36270 23580 36340
rect 23620 36270 23680 36340
rect 23720 36270 23780 36340
rect 23820 36270 23880 36340
rect 23920 36270 23980 36340
rect 24020 36270 24080 36340
rect 24120 36270 24180 36340
rect 24220 36270 24280 36340
rect 24320 36270 24380 36340
rect 24420 36270 24480 36340
rect 24520 36270 24580 36340
rect 24620 36270 24680 36340
rect 24720 36270 24780 36340
rect 24820 36270 24880 36340
rect 15200 36050 15300 36110
rect 6380 33980 6440 34040
rect 6480 33980 6540 34040
rect 6580 33980 6640 34040
rect 6680 33980 6740 34040
rect 6780 33980 6840 34040
rect 6880 33980 6940 34040
rect 6980 33980 7040 34040
rect 7080 33980 7140 34040
rect 7180 33980 7240 34040
rect 7280 33980 7340 34040
rect 7380 33980 7440 34040
rect 7480 33980 7540 34040
rect 7580 33980 7640 34040
rect 7680 33980 7740 34040
rect 7780 33980 7840 34040
rect 7880 33980 7940 34040
rect 7980 33980 8040 34040
rect 8080 33980 8140 34040
rect 8180 33980 8240 34040
rect 8280 33980 8340 34040
rect 8380 33980 8440 34040
rect 8480 33980 8540 34040
rect 8580 33980 8640 34040
rect 8680 33980 8740 34040
rect 8780 33980 8840 34040
rect 8880 33980 8940 34040
rect 8980 33980 9040 34040
rect 9080 33980 9140 34040
rect 9180 33980 9240 34040
rect 9280 33980 9340 34040
rect 9380 33980 9440 34040
rect 9480 33980 9540 34040
rect 9580 33980 9640 34040
rect 9680 33980 9740 34040
rect 9780 33980 9840 34040
rect 9880 33980 9940 34040
rect 9980 33980 10040 34040
rect 10080 33980 10140 34040
rect 10180 33980 10240 34040
rect 10280 33980 10340 34040
rect 10380 33980 10440 34040
rect 10480 33980 10540 34040
rect 10580 33980 10640 34040
rect 10680 33980 10740 34040
rect 10780 33980 10840 34040
rect 3810 33560 3870 33620
rect 3910 33560 3970 33620
rect 4010 33560 4070 33620
rect 4110 33560 4170 33620
rect 4210 33560 4270 33620
rect 4310 33560 4370 33620
rect 4410 33560 4470 33620
rect 4510 33560 4570 33620
rect 4610 33560 4670 33620
rect 4710 33560 4770 33620
rect 4810 33560 4870 33620
rect 4910 33560 4970 33620
rect 5010 33560 5070 33620
rect 5110 33560 5170 33620
rect 5210 33560 5270 33620
rect 5310 33560 5370 33620
rect 5410 33560 5470 33620
rect 5510 33560 5570 33620
rect 5610 33560 5670 33620
rect 5710 33560 5770 33620
rect 5810 33560 5870 33620
rect 5910 33560 5970 33620
rect 6010 33560 6070 33620
rect 6110 33560 6170 33620
rect 13768 32420 13848 32460
rect 16120 32110 16180 32180
rect 16220 32110 16280 32180
rect 16320 32110 16380 32180
rect 16420 32110 16480 32180
rect 16520 32110 16580 32180
rect 16620 32110 16680 32180
rect 16720 32110 16780 32180
rect 16820 32110 16880 32180
rect 16920 32110 16980 32180
rect 17020 32110 17080 32180
rect 17120 32110 17180 32180
rect 17220 32110 17280 32180
rect 17320 32110 17380 32180
rect 17420 32110 17480 32180
rect 17520 32110 17580 32180
rect 17620 32110 17680 32180
rect 17720 32110 17780 32180
rect 17820 32110 17880 32180
rect 17920 32110 17980 32180
rect 18020 32110 18080 32180
rect 18120 32110 18180 32180
rect 18220 32110 18280 32180
rect 18320 32110 18380 32180
rect 18420 32110 18480 32180
rect 18520 32110 18580 32180
rect 18620 32110 18680 32180
rect 18720 32110 18780 32180
rect 18820 32110 18880 32180
rect 18920 32110 18980 32180
rect 19020 32110 19080 32180
rect 19120 32110 19180 32180
rect 19220 32110 19280 32180
rect 19320 32110 19380 32180
rect 19420 32110 19480 32180
rect 19520 32110 19580 32180
rect 19620 32110 19680 32180
rect 19720 32110 19780 32180
rect 19820 32110 19880 32180
rect 19920 32110 19980 32180
rect 20020 32110 20080 32180
rect 20120 32110 20180 32180
rect 20220 32110 20280 32180
rect 20320 32110 20380 32180
rect 20420 32110 20480 32180
rect 20520 32110 20580 32180
rect 20620 32110 20680 32180
rect 20720 32110 20780 32180
rect 20820 32110 20880 32180
rect 20920 32110 20980 32180
rect 21020 32110 21080 32180
rect 21120 32110 21180 32180
rect 21220 32110 21280 32180
rect 21320 32110 21380 32180
rect 21420 32110 21480 32180
rect 21520 32110 21580 32180
rect 21620 32110 21680 32180
rect 21720 32110 21780 32180
rect 21820 32110 21880 32180
rect 21920 32110 21980 32180
rect 22020 32110 22080 32180
rect 22120 32110 22180 32180
rect 22220 32110 22280 32180
rect 22320 32110 22380 32180
rect 22420 32110 22480 32180
rect 22520 32110 22580 32180
rect 22620 32110 22680 32180
rect 22720 32110 22780 32180
rect 22820 32110 22880 32180
rect 22920 32110 22980 32180
rect 23020 32110 23080 32180
rect 23120 32110 23180 32180
rect 23220 32110 23280 32180
rect 23320 32110 23380 32180
rect 23420 32110 23480 32180
rect 23520 32110 23580 32180
rect 23620 32110 23680 32180
rect 23720 32110 23780 32180
rect 23820 32110 23880 32180
rect 23920 32110 23980 32180
rect 24020 32110 24080 32180
rect 24120 32110 24180 32180
rect 24220 32110 24280 32180
rect 24320 32110 24380 32180
rect 24420 32110 24480 32180
rect 24520 32110 24580 32180
rect 24620 32110 24680 32180
rect 24720 32110 24780 32180
rect 24820 32110 24880 32180
rect 24920 32110 24980 32180
rect 25020 32110 25080 32180
rect 25120 32110 25180 32180
rect 25220 32110 25280 32180
rect 25320 32110 25380 32180
rect 6440 29840 6500 29900
rect 6540 29840 6600 29900
rect 6640 29840 6700 29900
rect 6740 29840 6800 29900
rect 6840 29840 6900 29900
rect 6940 29840 7000 29900
rect 7040 29840 7100 29900
rect 7140 29840 7200 29900
rect 7240 29840 7300 29900
rect 7340 29840 7400 29900
rect 7440 29840 7500 29900
rect 7540 29840 7600 29900
rect 7640 29840 7700 29900
rect 7740 29840 7800 29900
rect 7840 29840 7900 29900
rect 7940 29840 8000 29900
rect 8040 29840 8100 29900
rect 8140 29840 8200 29900
rect 8240 29840 8300 29900
rect 8340 29840 8400 29900
rect 8440 29840 8500 29900
rect 8540 29840 8600 29900
rect 8640 29840 8700 29900
rect 8740 29840 8800 29900
rect 8840 29840 8900 29900
rect 8940 29840 9000 29900
rect 9040 29840 9100 29900
rect 9140 29840 9200 29900
rect 9240 29840 9300 29900
rect 9340 29840 9400 29900
rect 9440 29840 9500 29900
rect 9540 29840 9600 29900
rect 9640 29840 9700 29900
rect 9740 29840 9800 29900
rect 9840 29840 9900 29900
rect 9940 29840 10000 29900
rect 10040 29840 10100 29900
rect 10140 29840 10200 29900
rect 10240 29840 10300 29900
rect 10340 29840 10400 29900
rect 10440 29840 10500 29900
rect 10540 29840 10600 29900
rect 10640 29840 10700 29900
rect 10740 29840 10800 29900
rect 10840 29840 10900 29900
rect 10940 29840 11000 29900
rect 11040 29840 11100 29900
rect 11140 29840 11200 29900
rect 2210 29310 2270 29370
rect 2310 29310 2370 29370
rect 2410 29310 2470 29370
rect 2510 29310 2570 29370
rect 2610 29310 2670 29370
rect 2710 29310 2770 29370
rect 2810 29310 2870 29370
rect 2910 29310 2970 29370
rect 3010 29310 3070 29370
rect 3110 29310 3170 29370
rect 3210 29310 3270 29370
rect 3310 29310 3370 29370
rect 3410 29310 3470 29370
rect 3510 29310 3570 29370
rect 3610 29310 3670 29370
rect 3710 29310 3770 29370
rect 3810 29310 3870 29370
rect 3910 29310 3970 29370
rect 4010 29310 4070 29370
rect 4110 29310 4170 29370
rect 4210 29310 4270 29370
rect 4310 29310 4370 29370
rect 4410 29310 4470 29370
rect 4510 29310 4570 29370
rect 4610 29310 4670 29370
rect 4710 29310 4770 29370
rect 4810 29310 4870 29370
rect 4910 29310 4970 29370
rect 5010 29310 5070 29370
rect 5110 29310 5170 29370
rect 5210 29310 5270 29370
rect 5310 29310 5370 29370
rect 5410 29310 5470 29370
rect 5510 29310 5570 29370
rect 5610 29310 5670 29370
rect 5710 29310 5770 29370
rect 5810 29310 5870 29370
rect 5910 29310 5970 29370
rect 6010 29310 6070 29370
rect 6110 29310 6170 29370
rect 6210 29310 6270 29370
rect 7360 26570 7400 26610
rect 7440 26570 7480 26610
rect 7520 26570 7560 26610
rect 7600 26570 7640 26610
rect 7680 26570 7720 26610
rect 7760 26570 7800 26610
rect 7840 26570 7880 26610
rect 7920 26570 7960 26610
rect 8000 26570 8040 26610
rect 8080 26570 8120 26610
rect 8160 26570 8200 26610
rect 8240 26570 8280 26610
rect 8320 26570 8360 26610
rect 8400 26570 8440 26610
rect 8480 26570 8520 26610
rect 8560 26570 8600 26610
rect 8640 26570 8680 26610
rect 8720 26570 8760 26610
rect 8800 26570 8840 26610
rect 8880 26570 8920 26610
rect 8960 26570 9000 26610
rect 9040 26570 9080 26610
rect 9120 26570 9160 26610
rect 9200 26570 9240 26610
rect 9280 26570 9320 26610
rect 9360 26570 9400 26610
rect 9440 26570 9480 26610
rect 9520 26570 9560 26610
rect 9600 26570 9640 26610
rect 9680 26570 9720 26610
rect 9760 26570 9800 26610
rect 9840 26570 9880 26610
rect 9920 26570 9960 26610
rect 10000 26570 10040 26610
rect 10080 26570 10120 26610
rect 10160 26570 10200 26610
rect 10240 26570 10280 26610
rect 10320 26570 10360 26610
rect 10400 26570 10440 26610
rect 10480 26570 10520 26610
rect 10560 26570 10600 26610
rect 10640 26570 10680 26610
rect 10720 26570 10760 26610
rect 10800 26570 10840 26610
rect 10880 26570 10920 26610
rect 10960 26570 11000 26610
rect 11040 26570 11080 26610
rect 11120 26570 11160 26610
rect 11200 26570 11240 26610
rect 11280 26570 11320 26610
rect 11360 26570 11400 26610
rect 11440 26570 11480 26610
rect 11520 26570 11560 26610
rect 11600 26570 11640 26610
rect 11680 26570 11720 26610
rect 11760 26570 11800 26610
rect 11840 26570 11880 26610
rect 11920 26570 11960 26610
rect 12000 26570 12040 26610
rect 12080 26570 12120 26610
rect 12160 26570 12200 26610
rect 12240 26570 12280 26610
rect 12320 26570 12360 26610
rect 12400 26570 12440 26610
rect 12480 26570 12520 26610
rect 12560 26570 12600 26610
rect 12640 26570 12680 26610
rect 12720 26570 12760 26610
rect 12800 26570 12840 26610
rect 12880 26570 12920 26610
rect 12960 26570 13000 26610
rect 13040 26570 13080 26610
rect 13120 26570 13160 26610
rect 13200 26570 13240 26610
rect 13280 26570 13320 26610
rect 13360 26570 13400 26610
rect 13440 26570 13480 26610
rect 13520 26570 13560 26610
rect 13600 26570 13640 26610
rect 13680 26570 13720 26610
rect 13760 26570 13800 26610
rect 13840 26570 13880 26610
rect 13920 26570 13960 26610
rect 14000 26570 14040 26610
rect 14080 26570 14120 26610
rect 14160 26570 14200 26610
rect 14240 26570 14280 26610
rect 14320 26570 14360 26610
rect 14400 26570 14440 26610
rect 14480 26570 14520 26610
rect 14560 26570 14600 26610
rect 14640 26570 14680 26610
rect 14720 26570 14760 26610
rect 14800 26570 14840 26610
rect 14880 26570 14920 26610
rect 14960 26570 15000 26610
rect 15040 26570 15080 26610
rect 15120 26570 15160 26610
rect 15200 26570 15240 26610
rect 15280 26570 15320 26610
rect 15360 26570 15400 26610
rect 15440 26570 15480 26610
rect 15520 26570 15560 26610
rect 15600 26570 15640 26610
rect 15680 26570 15720 26610
rect 15760 26570 15800 26610
rect 15840 26570 15880 26610
rect 15920 26570 15960 26610
rect 16000 26570 16040 26610
rect 16080 26570 16120 26610
rect 16160 26570 16200 26610
rect 16240 26570 16280 26610
rect 16320 26570 16360 26610
rect 16400 26570 16440 26610
rect 16480 26570 16520 26610
rect 16560 26570 16600 26610
rect 16640 26570 16680 26610
rect 16720 26570 16760 26610
rect 16800 26570 16840 26610
rect 16880 26570 16920 26610
rect 16960 26570 17000 26610
rect 17040 26570 17080 26610
rect 17120 26570 17160 26610
rect 17200 26570 17240 26610
rect 17280 26570 17320 26610
rect 17360 26570 17400 26610
rect 17440 26570 17480 26610
rect 17520 26570 17560 26610
rect 17600 26570 17640 26610
rect 17680 26570 17720 26610
rect 17760 26570 17800 26610
rect 17840 26570 17880 26610
rect 17920 26570 17960 26610
rect 18000 26570 18040 26610
rect 18080 26570 18120 26610
rect 18160 26570 18200 26610
rect 18240 26570 18280 26610
rect 18320 26570 18360 26610
rect 18400 26570 18440 26610
rect 18480 26570 18520 26610
rect 18560 26570 18600 26610
rect 18640 26570 18680 26610
rect 18720 26570 18760 26610
rect 18800 26570 18840 26610
rect 18880 26570 18920 26610
rect 18960 26570 19000 26610
rect 19040 26570 19080 26610
rect 19120 26570 19160 26610
rect 19200 26570 19240 26610
rect 19280 26570 19320 26610
rect 19360 26570 19400 26610
rect 19440 26570 19480 26610
rect 19520 26570 19560 26610
rect 19600 26570 19640 26610
rect 19680 26570 19720 26610
rect 19760 26570 19800 26610
rect 19840 26570 19880 26610
rect 19920 26570 19960 26610
rect 20000 26570 20040 26610
rect 20080 26570 20120 26610
rect 20160 26570 20200 26610
rect 20240 26570 20280 26610
rect 20320 26570 20360 26610
rect 20400 26570 20440 26610
rect 20480 26570 20520 26610
rect 20560 26570 20600 26610
rect 7320 20960 7360 21000
rect 7400 20960 7440 21000
rect 7480 20960 7520 21000
rect 7560 20960 7600 21000
rect 7640 20960 7680 21000
rect 7720 20960 7760 21000
rect 7800 20960 7840 21000
rect 7880 20960 7920 21000
rect 7960 20960 8000 21000
rect 8040 20960 8080 21000
rect 8120 20960 8160 21000
rect 8200 20960 8240 21000
rect 8280 20960 8320 21000
rect 8360 20960 8400 21000
rect 8440 20960 8480 21000
rect 8520 20960 8560 21000
rect 8600 20960 8640 21000
rect 8680 20960 8720 21000
rect 8760 20960 8800 21000
rect 8840 20960 8880 21000
rect 8920 20960 8960 21000
rect 9000 20960 9040 21000
rect 9080 20960 9120 21000
rect 9160 20960 9200 21000
rect 9260 20960 9300 21000
rect 9340 20960 9380 21000
rect 9420 20960 9460 21000
rect 9500 20960 9540 21000
rect 9580 20960 9620 21000
rect 9660 20960 9700 21000
rect 9740 20960 9780 21000
rect 9820 20960 9860 21000
rect 9900 20960 9940 21000
rect 9980 20960 10020 21000
rect 10060 20960 10100 21000
rect 10140 20960 10180 21000
rect 10220 20960 10260 21000
rect 10300 20960 10340 21000
rect 10380 20960 10420 21000
rect 10460 20960 10500 21000
rect 10540 20960 10580 21000
rect 10620 20960 10660 21000
rect 10700 20960 10740 21000
rect 10780 20960 10820 21000
rect 10860 20960 10900 21000
rect 10940 20960 10980 21000
rect 11020 20960 11060 21000
rect 11100 20960 11140 21000
rect 11180 20960 11220 21000
rect 11260 20960 11300 21000
rect 11340 20960 11380 21000
rect 11420 20960 11460 21000
rect 11500 20960 11540 21000
rect 11580 20960 11620 21000
rect 11660 20960 11700 21000
rect 11740 20960 11780 21000
rect 11820 20960 11860 21000
rect 11900 20960 11940 21000
rect 11980 20960 12020 21000
rect 12060 20960 12100 21000
rect 12140 20960 12180 21000
rect 12220 20960 12260 21000
rect 12300 20960 12340 21000
rect 12380 20960 12420 21000
rect 12460 20960 12500 21000
rect 12540 20960 12580 21000
rect 12620 20960 12660 21000
rect 12700 20960 12740 21000
rect 12780 20960 12820 21000
rect 12880 20960 12920 21000
rect 12960 20960 13000 21000
rect 13040 20960 13080 21000
rect 13120 20960 13160 21000
rect 13200 20960 13240 21000
rect 13280 20960 13320 21000
rect 13360 20960 13400 21000
rect 13440 20960 13480 21000
rect 13520 20960 13560 21000
rect 13600 20960 13640 21000
rect 13680 20960 13720 21000
rect 13760 20960 13800 21000
rect 13840 20960 13880 21000
rect 13920 20960 13960 21000
rect 14000 20960 14040 21000
rect 14080 20960 14120 21000
rect 14160 20960 14200 21000
rect 14240 20960 14280 21000
rect 14320 20960 14360 21000
rect 14400 20960 14440 21000
rect 14480 20960 14520 21000
rect 14560 20960 14600 21000
rect 14640 20960 14680 21000
rect 14720 20960 14760 21000
rect 14800 20960 14840 21000
rect 14880 20960 14920 21000
rect 14960 20960 15000 21000
rect 15040 20960 15080 21000
rect 15120 20960 15160 21000
rect 15200 20960 15240 21000
rect 15280 20960 15320 21000
rect 15360 20960 15400 21000
rect 15440 20960 15480 21000
rect 15520 20960 15560 21000
rect 15600 20960 15640 21000
rect 15680 20960 15720 21000
rect 15760 20960 15800 21000
rect 15840 20960 15880 21000
rect 15920 20960 15960 21000
rect 16000 20960 16040 21000
rect 16080 20960 16120 21000
rect 16160 20960 16200 21000
rect 16240 20960 16280 21000
rect 16320 20960 16360 21000
rect 16400 20960 16440 21000
rect 16480 20960 16520 21000
rect 16560 20960 16600 21000
rect 16640 20960 16680 21000
rect 16720 20960 16760 21000
rect 16800 20960 16840 21000
rect 16880 20960 16920 21000
rect 16960 20960 17000 21000
rect 17040 20960 17080 21000
rect 17120 20960 17160 21000
rect 17200 20960 17240 21000
rect 17280 20960 17320 21000
rect 17360 20960 17400 21000
rect 17440 20960 17480 21000
rect 17520 20960 17560 21000
rect 17600 20960 17640 21000
rect 17680 20960 17720 21000
rect 17760 20960 17800 21000
rect 17840 20960 17880 21000
rect 17920 20960 17960 21000
rect 18000 20960 18040 21000
rect 18080 20960 18120 21000
rect 18160 20960 18200 21000
rect 18240 20960 18280 21000
rect 18320 20960 18360 21000
rect 18400 20960 18440 21000
rect 18480 20960 18520 21000
rect 18560 20960 18600 21000
rect 18640 20960 18680 21000
rect 18720 20960 18760 21000
rect 18800 20960 18840 21000
rect 18880 20960 18920 21000
rect 18960 20960 19000 21000
rect 19040 20960 19080 21000
rect 19120 20960 19160 21000
rect 19200 20960 19240 21000
rect 19280 20960 19320 21000
rect 19360 20960 19400 21000
rect 19440 20960 19480 21000
rect 19520 20960 19560 21000
rect 19600 20960 19640 21000
rect 19680 20960 19720 21000
rect 19760 20960 19800 21000
rect 19840 20960 19880 21000
rect 19920 20960 19960 21000
rect 20000 20960 20040 21000
rect 20080 20960 20120 21000
rect 20160 20960 20200 21000
rect 20240 20960 20280 21000
rect 20320 20960 20360 21000
rect 20400 20960 20440 21000
rect 20480 20960 20520 21000
rect 20560 20960 20600 21000
rect 7320 20430 7360 20470
rect 7400 20430 7440 20470
rect 7480 20430 7520 20470
rect 7560 20430 7600 20470
rect 7640 20430 7680 20470
rect 7720 20430 7760 20470
rect 7800 20430 7840 20470
rect 7880 20430 7920 20470
rect 7960 20430 8000 20470
rect 8040 20430 8080 20470
rect 8120 20430 8160 20470
rect 8360 19980 8400 20020
rect 8440 19980 8480 20020
rect 8520 19980 8560 20020
rect 8600 19980 8640 20020
rect 8680 19980 8720 20020
rect 8760 19980 8800 20020
rect 8840 19980 8880 20020
rect 8920 19980 8960 20020
rect 9000 19980 9040 20020
rect 9080 19980 9120 20020
rect 9160 19980 9200 20020
rect 9260 19980 9300 20020
rect 9340 19980 9380 20020
rect 9420 19980 9460 20020
rect 9500 19980 9540 20020
rect 9580 19980 9620 20020
rect 9660 19980 9700 20020
rect 9740 19980 9780 20020
rect 9820 19980 9860 20020
rect 9900 19980 9940 20020
rect 9980 19980 10020 20020
rect 10060 19980 10100 20020
rect 10140 19980 10180 20020
rect 10220 19980 10260 20020
rect 10300 19980 10340 20020
rect 10380 19980 10420 20020
rect 10460 19980 10500 20020
rect 10540 19980 10580 20020
rect 10620 19980 10660 20020
rect 10700 19980 10740 20020
rect 10780 19980 10820 20020
rect 10860 19980 10900 20020
rect 10940 19980 10980 20020
rect 11020 19980 11060 20020
rect 11100 19980 11140 20020
rect 11180 19980 11220 20020
rect 11260 19980 11300 20020
rect 11340 19980 11380 20020
rect 11420 19980 11460 20020
rect 11500 19980 11540 20020
rect 11580 19980 11620 20020
rect 11660 19980 11700 20020
rect 11740 19980 11780 20020
rect 11820 19980 11860 20020
rect 11900 19980 11940 20020
rect 11980 19980 12020 20020
rect 12060 19980 12100 20020
rect 12140 19980 12180 20020
rect 12220 19980 12260 20020
rect 12300 19980 12340 20020
rect 12380 19980 12420 20020
rect 12460 19980 12500 20020
rect 12540 19980 12580 20020
rect 12620 19980 12660 20020
rect 12700 19980 12740 20020
rect 12780 19980 12820 20020
rect 12860 19980 12900 20020
rect 12940 19980 12980 20020
rect 13040 19980 13080 20020
rect 13120 19980 13160 20020
rect 13200 19980 13240 20020
rect 13280 19980 13320 20020
rect 13360 19980 13400 20020
rect 13440 19980 13480 20020
rect 13520 19980 13560 20020
rect 13600 19980 13640 20020
rect 13680 19980 13720 20020
rect 13760 19980 13800 20020
rect 13840 19980 13880 20020
rect 13920 19980 13960 20020
rect 14000 19980 14040 20020
rect 14080 19980 14120 20020
rect 14160 19980 14200 20020
rect 14240 19980 14280 20020
rect 14320 19980 14360 20020
rect 14400 19980 14440 20020
rect 14480 19980 14520 20020
rect 14560 19980 14600 20020
rect 14640 19980 14680 20020
rect 14720 19980 14760 20020
rect 14800 19980 14840 20020
rect 14880 19980 14920 20020
rect 14960 19980 15000 20020
rect 15040 19980 15080 20020
rect 15120 19980 15160 20020
rect 15200 19980 15240 20020
rect 15280 19980 15320 20020
rect 15360 19980 15400 20020
rect 15440 19980 15480 20020
rect 15520 19980 15560 20020
rect 15600 19980 15640 20020
rect 15680 19980 15720 20020
rect 15760 19980 15800 20020
rect 15840 19980 15880 20020
rect 15920 19980 15960 20020
rect 16000 19980 16040 20020
rect 16080 19980 16120 20020
rect 16160 19980 16200 20020
rect 16240 19980 16280 20020
rect 16320 19980 16360 20020
rect 16400 19980 16440 20020
rect 16480 19980 16520 20020
rect 16560 19980 16600 20020
rect 16640 19980 16680 20020
rect 16720 19980 16760 20020
rect 16800 19980 16840 20020
rect 16880 19980 16920 20020
rect 16960 19980 17000 20020
rect 17040 19980 17080 20020
rect 17120 19980 17160 20020
rect 17200 19980 17240 20020
rect 17280 19980 17320 20020
rect 17360 19980 17400 20020
rect 17440 19980 17480 20020
rect 17520 19980 17560 20020
rect 17600 19980 17640 20020
rect 17680 19980 17720 20020
rect 17760 19980 17800 20020
rect 17840 19980 17880 20020
rect 17920 19980 17960 20020
rect 18000 19980 18040 20020
rect 18080 19980 18120 20020
rect 18160 19980 18200 20020
rect 18240 19980 18280 20020
rect 18320 19980 18360 20020
rect 18400 19980 18440 20020
rect 18480 19980 18520 20020
rect 18560 19980 18600 20020
rect 18640 19980 18680 20020
rect 18720 19980 18760 20020
rect 18800 19980 18840 20020
rect 18880 19980 18920 20020
rect 18960 19980 19000 20020
rect 19040 19980 19080 20020
rect 19120 19980 19160 20020
rect 19200 19980 19240 20020
rect 19280 19980 19320 20020
rect 19360 19980 19400 20020
rect 19440 19980 19480 20020
rect 19520 19980 19560 20020
rect 19600 19980 19640 20020
rect 19680 19980 19720 20020
rect 19760 19980 19800 20020
rect 19840 19980 19880 20020
rect 19920 19980 19960 20020
rect 20000 19980 20040 20020
rect 20080 19980 20120 20020
rect 20160 19980 20200 20020
rect 20240 19980 20280 20020
rect 20320 19980 20360 20020
rect 20400 19980 20440 20020
rect 20480 19980 20520 20020
rect 20560 19980 20600 20020
rect 9700 14300 9740 14340
rect 9790 14300 9830 14340
rect 9870 14300 9910 14340
rect 9950 14300 9990 14340
rect 10030 14300 10070 14340
rect 10110 14300 10150 14340
rect 10190 14300 10230 14340
rect 10270 14300 10310 14340
rect 10350 14300 10390 14340
rect 10430 14300 10470 14340
rect 10510 14300 10550 14340
rect 10590 14300 10630 14340
rect 10670 14300 10710 14340
rect 10750 14300 10790 14340
rect 10830 14300 10870 14340
rect 10910 14300 10950 14340
rect 10990 14300 11030 14340
rect 11070 14300 11110 14340
rect 11150 14300 11190 14340
rect 11230 14300 11270 14340
rect 11310 14300 11350 14340
rect 11390 14300 11430 14340
rect 11470 14300 11510 14340
rect 11550 14300 11590 14340
rect 11630 14300 11670 14340
rect 11710 14300 11750 14340
rect 11790 14300 11830 14340
rect 11870 14300 11910 14340
rect 11950 14300 11990 14340
rect 12030 14300 12070 14340
rect 12110 14300 12150 14340
rect 12190 14300 12230 14340
rect 12270 14300 12310 14340
rect 12350 14300 12390 14340
rect 12430 14300 12470 14340
rect 12510 14300 12550 14340
rect 12590 14300 12630 14340
rect 12670 14300 12710 14340
rect 12750 14300 12790 14340
rect 12830 14300 12870 14340
rect 12910 14300 12950 14340
rect 12990 14300 13030 14340
rect 13070 14300 13110 14340
rect 13150 14300 13230 14340
rect 13270 14300 13310 14340
rect 13350 14300 13390 14340
rect 13430 14300 13470 14340
rect 13510 14300 13550 14340
rect 13590 14300 13630 14340
rect 13670 14300 13710 14340
rect 13750 14300 13790 14340
rect 13830 14300 13870 14340
rect 13910 14300 13950 14340
rect 13990 14300 14030 14340
rect 14070 14300 14110 14340
rect 14150 14300 14190 14340
rect 14230 14300 14270 14340
rect 14310 14300 14350 14340
rect 14390 14300 14430 14340
rect 14470 14300 14510 14340
rect 14550 14300 14590 14340
rect 14630 14300 14670 14340
rect 14710 14300 14750 14340
rect 14790 14300 14830 14340
rect 14870 14300 14910 14340
rect 14950 14300 14990 14340
rect 15030 14300 15070 14340
rect 15110 14300 15150 14340
rect 15190 14300 15230 14340
rect 15270 14300 15310 14340
rect 15350 14300 15390 14340
rect 15430 14300 15470 14340
rect 15510 14300 15550 14340
rect 15590 14300 15630 14340
rect 15670 14300 15710 14340
rect 15750 14300 15790 14340
rect 15830 14300 15870 14340
rect 15910 14300 15950 14340
rect 15990 14300 16030 14340
rect 16070 14300 16110 14340
rect 16150 14300 16190 14340
rect 16230 14300 16270 14340
rect 16310 14300 16350 14340
rect 16390 14300 16430 14340
rect 16470 14300 16510 14340
rect 16550 14300 16590 14340
rect 16630 14300 16670 14340
rect 16710 14300 16750 14340
rect 16790 14300 16830 14340
rect 16870 14300 16910 14340
rect 16950 14300 16990 14340
rect 17030 14300 17070 14340
rect 17110 14300 17150 14340
rect 17190 14300 17230 14340
rect 17270 14300 17310 14340
rect 17350 14300 17390 14340
rect 17430 14300 17470 14340
rect 17510 14300 17550 14340
rect 17590 14300 17630 14340
rect 17670 14300 17710 14340
rect 17750 14300 17790 14340
rect 17830 14300 17870 14340
rect 17910 14300 17950 14340
rect 17990 14300 18030 14340
rect 18070 14300 18110 14340
rect 18150 14300 18190 14340
rect 18230 14300 18270 14340
rect 18310 14300 18350 14340
rect 18390 14300 18430 14340
rect 18470 14300 18510 14340
rect 18550 14300 18590 14340
rect 18630 14300 18670 14340
rect 18710 14300 18750 14340
rect 18790 14300 18830 14340
rect 18870 14300 18910 14340
rect 18950 14300 18990 14340
rect 19030 14300 19070 14340
rect 19110 14300 19150 14340
rect 19190 14300 19230 14340
rect 19270 14300 19310 14340
rect 19350 14300 19390 14340
rect 19430 14300 19470 14340
rect 19510 14300 19550 14340
rect 19590 14300 19630 14340
rect 19670 14300 19710 14340
rect 19750 14300 19790 14340
rect 19830 14300 19870 14340
rect 19910 14300 19950 14340
rect 19990 14300 20030 14340
rect 20070 14300 20110 14340
rect 20150 14300 20190 14340
rect 20230 14300 20270 14340
rect 20310 14300 20350 14340
rect 20390 14300 20430 14340
rect 20470 14300 20510 14340
rect 20550 14300 20590 14340
rect 20630 14300 20670 14340
rect 20710 14300 20750 14340
rect 20790 14300 20830 14340
rect 20870 14300 20910 14340
rect 20950 14300 20990 14340
rect 21030 14300 21070 14340
rect 7320 13330 7360 13370
rect 7400 13330 7440 13370
rect 7480 13330 7520 13370
rect 7560 13330 7600 13370
rect 7640 13330 7680 13370
rect 7720 13330 7760 13370
rect 7800 13330 7840 13370
rect 7880 13330 7920 13370
rect 7960 13330 8000 13370
rect 8040 13330 8080 13370
rect 8120 13330 8160 13370
rect 8200 13330 8240 13370
rect 8280 13330 8320 13370
rect 8360 13330 8400 13370
rect 8440 13330 8480 13370
rect 8520 13330 8560 13370
rect 8600 13330 8640 13370
rect 8680 13330 8720 13370
rect 8760 13330 8800 13370
rect 8840 13330 8880 13370
rect 8920 13330 8960 13370
rect 9000 13330 9040 13370
rect 9080 13330 9120 13370
rect 9160 13330 9200 13370
rect 9240 13330 9280 13370
rect 9320 13330 9360 13370
rect 9400 13330 9440 13370
rect 9480 13330 9520 13370
rect 9560 13330 9600 13370
rect 9640 13330 9680 13370
rect 9720 13330 9760 13370
rect 9800 13330 9840 13370
rect 9890 13330 9930 13370
rect 9970 13330 10010 13370
rect 10050 13330 10090 13370
rect 10130 13330 10170 13370
rect 10210 13330 10250 13370
rect 10290 13330 10330 13370
rect 10370 13330 10410 13370
rect 10450 13330 10490 13370
rect 10530 13330 10570 13370
rect 10610 13330 10650 13370
rect 10690 13330 10730 13370
rect 10770 13330 10810 13370
rect 10850 13330 10890 13370
rect 10930 13330 10970 13370
rect 11010 13330 11050 13370
rect 11090 13330 11130 13370
rect 11170 13330 11210 13370
rect 11250 13330 11290 13370
rect 11330 13330 11370 13370
rect 11410 13330 11450 13370
rect 11490 13330 11530 13370
rect 11570 13330 11610 13370
rect 11650 13330 11690 13370
rect 11730 13330 11770 13370
rect 11810 13330 11850 13370
rect 11890 13330 11930 13370
rect 11970 13330 12010 13370
rect 12050 13330 12090 13370
rect 12130 13330 12170 13370
rect 12210 13330 12250 13370
rect 12290 13330 12330 13370
rect 12370 13330 12410 13370
rect 12450 13330 12490 13370
rect 12530 13330 12570 13370
rect 12610 13330 12650 13370
rect 12690 13330 12730 13370
rect 12770 13330 12810 13370
rect 12850 13330 12890 13370
rect 12930 13330 12970 13370
rect 13010 13330 13050 13370
rect 13090 13330 13130 13370
rect 13170 13330 13210 13370
rect 13250 13330 13290 13370
rect 13330 13330 13400 13370
rect 13440 13330 13480 13370
rect 13520 13330 13560 13370
rect 13600 13330 13640 13370
rect 13680 13330 13720 13370
rect 13760 13330 13800 13370
rect 13840 13330 13880 13370
rect 13920 13330 13960 13370
rect 14000 13330 14040 13370
rect 14080 13330 14120 13370
rect 14160 13330 14200 13370
rect 14240 13330 14280 13370
rect 14320 13330 14360 13370
rect 14400 13330 14440 13370
rect 14480 13330 14520 13370
rect 14560 13330 14600 13370
rect 14640 13330 14680 13370
rect 14720 13330 14760 13370
rect 14800 13330 14840 13370
rect 14880 13330 14920 13370
rect 14960 13330 15000 13370
rect 15040 13330 15080 13370
rect 15120 13330 15160 13370
rect 15200 13330 15240 13370
rect 15280 13330 15320 13370
rect 15360 13330 15400 13370
rect 15440 13330 15480 13370
rect 15520 13330 15560 13370
rect 15600 13330 15640 13370
rect 15680 13330 15720 13370
rect 15760 13330 15800 13370
rect 15840 13330 15880 13370
rect 15920 13330 15960 13370
rect 16000 13330 16040 13370
rect 16080 13330 16120 13370
rect 16160 13330 16200 13370
rect 16240 13330 16280 13370
rect 16320 13330 16360 13370
rect 16400 13330 16440 13370
rect 16480 13330 16520 13370
rect 16560 13330 16600 13370
rect 16640 13330 16680 13370
rect 16720 13330 16760 13370
rect 16800 13330 16840 13370
rect 16880 13330 16920 13370
rect 16960 13330 17000 13370
rect 17040 13330 17080 13370
rect 17120 13330 17160 13370
rect 17200 13330 17240 13370
rect 17280 13330 17320 13370
rect 17360 13330 17400 13370
rect 17440 13330 17480 13370
rect 17520 13330 17560 13370
rect 17600 13330 17640 13370
rect 17680 13330 17720 13370
rect 17760 13330 17800 13370
rect 17840 13330 17880 13370
rect 17920 13330 17960 13370
rect 18000 13330 18040 13370
rect 18080 13330 18120 13370
rect 18160 13330 18200 13370
rect 18240 13330 18280 13370
rect 18320 13330 18360 13370
rect 18400 13330 18440 13370
rect 18480 13330 18520 13370
rect 18560 13330 18600 13370
rect 18640 13330 18680 13370
rect 18720 13330 18760 13370
rect 18800 13330 18840 13370
rect 18880 13330 18920 13370
rect 18960 13330 19000 13370
rect 19040 13330 19080 13370
rect 19120 13330 19160 13370
rect 19200 13330 19240 13370
rect 19280 13330 19320 13370
rect 19360 13330 19400 13370
rect 19440 13330 19480 13370
rect 19520 13330 19560 13370
rect 19600 13330 19640 13370
rect 19680 13330 19720 13370
rect 19760 13330 19800 13370
rect 19840 13330 19880 13370
rect 19920 13330 19960 13370
rect 20000 13330 20040 13370
rect 20080 13330 20120 13370
rect 20160 13330 20200 13370
rect 20240 13330 20280 13370
rect 20320 13330 20360 13370
rect 20400 13330 20440 13370
rect 20480 13330 20520 13370
rect 20560 13330 20600 13370
rect 20640 13330 20680 13370
rect 20720 13330 20760 13370
rect 20800 13330 20840 13370
rect 20880 13330 20920 13370
rect 20960 13330 21000 13370
rect 21040 13330 21080 13370
rect 7320 9680 7360 9720
rect 7400 9680 7440 9720
rect 7480 9680 7520 9720
rect 7560 9680 7600 9720
rect 7640 9680 7680 9720
rect 7720 9680 7760 9720
rect 8520 9680 8560 9720
rect 8600 9680 8640 9720
rect 8680 9680 8720 9720
rect 8760 9680 8800 9720
rect 8840 9680 8880 9720
rect 8920 9680 8960 9720
rect 9000 9680 9040 9720
rect 9080 9680 9120 9720
rect 9160 9680 9200 9720
rect 9240 9680 9280 9720
rect 9320 9680 9360 9720
rect 9400 9680 9440 9720
rect 9480 9680 9520 9720
rect 9560 9680 9600 9720
rect 9640 9680 9680 9720
rect 9720 9680 9760 9720
rect 9800 9680 9840 9720
rect 9890 9680 9930 9720
rect 9970 9680 10010 9720
rect 10050 9680 10090 9720
rect 10130 9680 10170 9720
rect 10210 9680 10250 9720
rect 10290 9680 10330 9720
rect 10370 9680 10410 9720
rect 10450 9680 10490 9720
rect 10530 9680 10570 9720
rect 10610 9680 10650 9720
rect 10690 9680 10730 9720
rect 10770 9680 10810 9720
rect 10850 9680 10890 9720
rect 10930 9680 10970 9720
rect 11010 9680 11050 9720
rect 11090 9680 11130 9720
rect 11170 9680 11210 9720
rect 11250 9680 11290 9720
rect 11330 9680 11370 9720
rect 11410 9680 11450 9720
rect 11490 9680 11530 9720
rect 11570 9680 11610 9720
rect 11650 9680 11690 9720
rect 11730 9680 11770 9720
rect 11810 9680 11850 9720
rect 11890 9680 11930 9720
rect 11970 9680 12010 9720
rect 12050 9680 12090 9720
rect 12130 9680 12170 9720
rect 12210 9680 12250 9720
rect 12290 9680 12330 9720
rect 12370 9680 12410 9720
rect 12450 9680 12490 9720
rect 12530 9680 12570 9720
rect 12610 9680 12650 9720
rect 12690 9680 12730 9720
rect 12770 9680 12810 9720
rect 12850 9680 12890 9720
rect 12930 9680 12970 9720
rect 13010 9680 13050 9720
rect 13090 9680 13130 9720
rect 13170 9680 13210 9720
rect 13250 9680 13290 9720
rect 13330 9680 13370 9720
rect 13410 9680 13450 9720
rect 13490 9680 13530 9720
rect 13570 9680 13610 9720
rect 13650 9680 13690 9720
rect 13730 9680 13770 9720
rect 13810 9680 13850 9720
rect 13890 9680 13930 9720
rect 13970 9680 14010 9720
rect 14050 9680 14090 9720
rect 14130 9680 14170 9720
rect 14210 9680 14250 9720
rect 14290 9680 14330 9720
rect 14370 9680 14410 9720
rect 14450 9680 14490 9720
rect 14530 9680 14570 9720
rect 14610 9680 14650 9720
rect 14690 9680 14730 9720
rect 14770 9680 14810 9720
rect 14850 9680 14890 9720
rect 14930 9680 14970 9720
rect 15010 9680 15050 9720
rect 15090 9680 15130 9720
rect 15170 9680 15210 9720
rect 15250 9680 15290 9720
rect 15330 9680 15370 9720
rect 15410 9680 15450 9720
rect 15490 9680 15530 9720
rect 15570 9680 15610 9720
rect 15650 9680 15690 9720
rect 15730 9680 15770 9720
rect 15810 9680 15850 9720
rect 15890 9680 15930 9720
rect 15970 9680 16010 9720
rect 16050 9680 16090 9720
rect 16130 9680 16170 9720
rect 16210 9680 16250 9720
rect 16290 9680 16330 9720
rect 16370 9680 16410 9720
rect 16450 9680 16490 9720
rect 16530 9680 16570 9720
rect 16610 9680 16650 9720
rect 16690 9680 16730 9720
rect 16770 9680 16810 9720
rect 16850 9680 16890 9720
rect 16930 9680 16970 9720
rect 17010 9680 17050 9720
rect 17090 9680 17130 9720
rect 17170 9680 17210 9720
rect 17250 9680 17290 9720
rect 17330 9680 17370 9720
rect 17410 9680 17450 9720
rect 17490 9680 17530 9720
rect 17570 9680 17610 9720
rect 17650 9680 17690 9720
rect 17730 9680 17770 9720
rect 17810 9680 17850 9720
rect 17890 9680 17930 9720
rect 17970 9680 18010 9720
rect 18050 9680 18090 9720
rect 18130 9680 18170 9720
rect 18210 9680 18250 9720
rect 18290 9680 18330 9720
rect 18370 9680 18410 9720
rect 18450 9680 18490 9720
rect 18530 9680 18570 9720
rect 18610 9680 18650 9720
rect 18690 9680 18730 9720
rect 18770 9680 18810 9720
rect 18850 9680 18890 9720
rect 18930 9680 18970 9720
rect 19010 9680 19050 9720
rect 19090 9680 19130 9720
rect 19170 9680 19210 9720
rect 19250 9680 19290 9720
rect 19330 9680 19370 9720
rect 19410 9680 19450 9720
rect 19490 9680 19530 9720
rect 19570 9680 19610 9720
rect 19650 9680 19690 9720
rect 19730 9680 19770 9720
rect 19810 9680 19850 9720
rect 19890 9680 19930 9720
rect 19970 9680 20010 9720
rect 20050 9680 20090 9720
rect 20130 9680 20170 9720
rect 20210 9680 20250 9720
rect 20290 9680 20330 9720
rect 20370 9680 20410 9720
rect 20450 9680 20490 9720
rect 20530 9680 20570 9720
rect 20610 9680 20650 9720
rect 20690 9680 20730 9720
rect 20770 9680 20810 9720
rect 20850 9680 20890 9720
rect 20930 9680 20970 9720
rect 21010 9680 21050 9720
rect 7740 9590 7780 9630
rect 7820 9590 7860 9630
rect 7900 9590 7940 9630
rect 7980 9590 8020 9630
rect 8060 9590 8100 9630
rect 8140 9590 8180 9630
rect 8220 9590 8260 9630
rect 8300 9590 8340 9630
rect 8380 9590 8420 9630
rect 8460 9590 8500 9630
rect 9900 6930 9960 6980
rect 10120 6930 10180 6980
rect 10340 6930 10400 6980
rect 10560 6930 10620 6980
rect 10780 6930 10840 6980
rect 11000 6930 11060 6980
rect 11220 6930 11280 6980
rect 11440 6930 11500 6980
rect 11660 6930 11720 6980
rect 11880 6930 11940 6980
rect 12100 6930 12160 6980
rect 12320 6930 12380 6980
rect 12540 6930 12600 6980
rect 12760 6930 12820 6980
rect 12980 6930 13040 6980
rect 13200 6930 13260 6980
rect 13670 6930 13730 6980
rect 13890 6930 13950 6980
rect 14110 6930 14170 6980
rect 14330 6930 14390 6980
rect 14550 6930 14610 6980
rect 14770 6930 14830 6980
rect 14990 6930 15050 6980
rect 15210 6930 15270 6980
rect 15430 6930 15490 6980
rect 15650 6930 15710 6980
rect 15870 6930 15930 6980
rect 16090 6930 16150 6980
rect 16310 6930 16370 6980
rect 16530 6930 16590 6980
rect 16750 6930 16810 6980
rect 16970 6930 17030 6980
rect 13630 5940 13690 5990
rect 13850 5940 13910 5990
rect 14070 5940 14130 5990
rect 14290 5940 14350 5990
rect 14510 5940 14570 5990
rect 14730 5940 14790 5990
rect 14950 5940 15010 5990
rect 15170 5940 15230 5990
rect 15390 5940 15450 5990
rect 15610 5940 15670 5990
rect 15830 5940 15890 5990
rect 16050 5940 16110 5990
rect 16270 5940 16330 5990
rect 16490 5940 16550 5990
rect 16710 5940 16770 5990
rect 16930 5940 16990 5990
rect 9930 5830 9970 5870
rect 10010 5830 10050 5870
rect 10090 5830 10130 5870
rect 10170 5830 10210 5870
rect 10250 5830 10290 5870
rect 10330 5830 10370 5870
rect 10410 5830 10450 5870
rect 10490 5830 10530 5870
rect 10610 5830 10650 5870
rect 10690 5830 10730 5870
rect 10770 5830 10810 5870
rect 10850 5830 10890 5870
rect 10930 5830 10970 5870
rect 11010 5830 11050 5870
rect 11090 5830 11130 5870
rect 11170 5830 11210 5870
rect 11250 5830 11290 5870
rect 11370 5830 11410 5870
rect 11450 5830 11490 5870
rect 11530 5830 11570 5870
rect 11610 5830 11650 5870
rect 11690 5830 11730 5870
rect 11770 5830 11810 5870
rect 11850 5830 11890 5870
rect 11930 5830 11970 5870
rect 12010 5830 12050 5870
rect 12130 5830 12170 5870
rect 12210 5830 12250 5870
rect 12290 5830 12330 5870
rect 12370 5830 12410 5870
rect 12450 5830 12490 5870
rect 12530 5830 12570 5870
rect 12610 5830 12650 5870
rect 12690 5830 12730 5870
rect 12770 5830 12810 5870
rect 12850 5830 12890 5870
rect 12930 5830 12970 5870
rect 13010 5830 13050 5870
rect 13090 5830 13130 5870
<< poly >>
rect 23530 43180 23560 43210
rect 21790 42880 21820 42910
rect 22020 42880 22050 42910
rect 22650 42890 22680 42920
rect 22950 42890 22980 42920
rect 23060 42890 23090 42920
rect 23530 42330 23560 42480
rect 23450 42320 23560 42330
rect 23450 42280 23470 42320
rect 23510 42280 23560 42320
rect 23450 42270 23560 42280
rect 23450 42210 23560 42220
rect 2739 42050 2849 42060
rect 2739 42010 2789 42050
rect 2829 42010 2849 42050
rect 2739 42000 2849 42010
rect 2629 41920 2659 41950
rect 2739 41920 2769 42000
rect 21790 41980 21820 42180
rect 22020 42140 22050 42180
rect 22020 42130 22150 42140
rect 22020 42080 22070 42130
rect 22050 42070 22070 42080
rect 22130 42070 22150 42130
rect 22650 42110 22680 42190
rect 22050 42060 22150 42070
rect 22570 42100 22680 42110
rect 22570 42060 22590 42100
rect 22630 42060 22680 42100
rect 22570 42050 22680 42060
rect 22950 42040 22980 42190
rect 23060 42150 23090 42190
rect 23450 42170 23500 42210
rect 23540 42170 23560 42210
rect 23450 42160 23560 42170
rect 23060 42140 23170 42150
rect 23060 42100 23110 42140
rect 23150 42100 23170 42140
rect 23450 42100 23480 42160
rect 23060 42090 23170 42100
rect 22950 42030 23060 42040
rect 22950 41990 23000 42030
rect 23040 41990 23060 42030
rect 22950 41980 23060 41990
rect 2849 41920 2879 41950
rect 21790 41970 21910 41980
rect 21790 41930 21850 41970
rect 21890 41930 21910 41970
rect 21790 41920 21910 41930
rect 21790 41880 21820 41920
rect 22950 41910 23060 41920
rect 3459 41820 3489 41850
rect 3569 41820 3599 41850
rect 3679 41820 3709 41850
rect 3789 41820 3819 41850
rect 3899 41820 3929 41850
rect 4009 41820 4039 41850
rect 4119 41820 4149 41850
rect 4229 41820 4259 41850
rect 6019 41840 6049 41870
rect 6249 41840 6279 41870
rect 6359 41840 6389 41870
rect 6589 41840 6619 41870
rect 6699 41840 6729 41870
rect 6809 41840 6839 41870
rect 6919 41840 6949 41870
rect 7149 41840 7179 41870
rect 7259 41840 7289 41870
rect 7369 41840 7399 41870
rect 7479 41840 7509 41870
rect 7589 41840 7619 41870
rect 7699 41840 7729 41870
rect 7809 41840 7839 41870
rect 7919 41840 7949 41870
rect 8209 41840 8239 41870
rect 8319 41840 8349 41870
rect 8429 41840 8459 41870
rect 8539 41840 8569 41870
rect 8649 41840 8679 41870
rect 8759 41840 8789 41870
rect 8869 41840 8899 41870
rect 8979 41840 9009 41870
rect 9089 41840 9119 41870
rect 9199 41840 9229 41870
rect 9309 41840 9339 41870
rect 9419 41840 9449 41870
rect 9529 41840 9559 41870
rect 9639 41840 9669 41870
rect 9749 41840 9779 41870
rect 9859 41840 9889 41870
rect 2629 41630 2659 41720
rect 2739 41690 2769 41720
rect 2629 41620 2739 41630
rect 2629 41580 2679 41620
rect 2719 41580 2739 41620
rect 2629 41570 2739 41580
rect 2849 41590 2879 41720
rect 2849 41580 2959 41590
rect 2849 41540 2899 41580
rect 2939 41540 2959 41580
rect 2849 41530 2959 41540
rect 2509 41400 2539 41430
rect 2619 41400 2649 41430
rect 2729 41400 2759 41430
rect 2839 41400 2869 41430
rect 2949 41400 2979 41430
rect 4609 41810 4639 41840
rect 4719 41810 4749 41840
rect 4829 41810 4859 41840
rect 4939 41810 4969 41840
rect 5049 41810 5079 41840
rect 5159 41810 5189 41840
rect 5269 41810 5299 41840
rect 5379 41810 5409 41840
rect 3459 41040 3489 41070
rect 3569 41040 3599 41070
rect 3679 41040 3709 41070
rect 3789 41040 3819 41070
rect 3899 41040 3929 41070
rect 4009 41040 4039 41070
rect 4119 41040 4149 41070
rect 4229 41040 4259 41070
rect 22950 41870 23000 41910
rect 23040 41870 23060 41910
rect 23450 41870 23480 41900
rect 22950 41860 23060 41870
rect 22570 41800 22680 41810
rect 22570 41760 22590 41800
rect 22630 41760 22680 41800
rect 22570 41750 22680 41760
rect 22650 41710 22680 41750
rect 22950 41710 22980 41860
rect 23060 41800 23170 41810
rect 23060 41760 23110 41800
rect 23150 41760 23170 41800
rect 23060 41750 23170 41760
rect 23450 41760 23560 41770
rect 23060 41710 23090 41750
rect 23450 41720 23500 41760
rect 23540 41720 23560 41760
rect 23450 41710 23560 41720
rect 21790 41650 21820 41680
rect 23450 41570 23480 41710
rect 22650 41480 22680 41510
rect 22950 41480 22980 41510
rect 23060 41480 23090 41510
rect 23450 41340 23480 41370
rect 6019 41300 6049 41340
rect 6249 41300 6279 41340
rect 5959 41280 6049 41300
rect 5959 41240 5969 41280
rect 6009 41240 6049 41280
rect 5959 41220 6049 41240
rect 6189 41280 6279 41300
rect 6189 41240 6199 41280
rect 6239 41260 6279 41280
rect 6359 41260 6389 41340
rect 6589 41300 6619 41340
rect 6239 41240 6389 41260
rect 6189 41220 6389 41240
rect 6529 41280 6619 41300
rect 6529 41240 6539 41280
rect 6579 41260 6619 41280
rect 6699 41260 6729 41340
rect 6809 41260 6839 41340
rect 6919 41260 6949 41340
rect 7149 41300 7179 41340
rect 6579 41240 6949 41260
rect 6529 41220 6949 41240
rect 7089 41280 7179 41300
rect 7089 41240 7099 41280
rect 7139 41260 7179 41280
rect 7259 41260 7289 41340
rect 7369 41260 7399 41340
rect 7479 41260 7509 41340
rect 7589 41260 7619 41340
rect 7699 41260 7729 41340
rect 7809 41260 7839 41340
rect 7919 41260 7949 41340
rect 8209 41300 8239 41340
rect 7139 41240 7949 41260
rect 7089 41220 7949 41240
rect 8149 41280 8239 41300
rect 8149 41240 8159 41280
rect 8199 41260 8239 41280
rect 8319 41260 8349 41340
rect 8429 41260 8459 41340
rect 8539 41260 8569 41340
rect 8649 41260 8679 41340
rect 8759 41260 8789 41340
rect 8869 41260 8899 41340
rect 8979 41260 9009 41340
rect 9089 41260 9119 41340
rect 9199 41260 9229 41340
rect 9309 41260 9339 41340
rect 9419 41260 9449 41340
rect 9529 41260 9559 41340
rect 9639 41260 9669 41340
rect 9749 41260 9779 41340
rect 9859 41260 9889 41340
rect 8199 41240 9889 41260
rect 8149 41220 9889 41240
rect 6019 41180 6049 41220
rect 6249 41180 6279 41220
rect 6359 41180 6389 41220
rect 6589 41180 6619 41220
rect 6699 41180 6729 41220
rect 6809 41180 6839 41220
rect 6919 41180 6949 41220
rect 7149 41180 7179 41220
rect 7259 41180 7289 41220
rect 7369 41180 7399 41220
rect 7479 41180 7509 41220
rect 7589 41180 7619 41220
rect 7699 41180 7729 41220
rect 7809 41180 7839 41220
rect 7919 41180 7949 41220
rect 8209 41180 8239 41220
rect 8319 41180 8349 41220
rect 8429 41180 8459 41220
rect 8539 41180 8569 41220
rect 8649 41180 8679 41220
rect 8759 41180 8789 41220
rect 8869 41180 8899 41220
rect 8979 41180 9009 41220
rect 9089 41180 9119 41220
rect 9199 41180 9229 41220
rect 9309 41180 9339 41220
rect 9419 41180 9449 41220
rect 9529 41180 9559 41220
rect 9639 41180 9669 41220
rect 9749 41180 9779 41220
rect 9859 41180 9889 41220
rect 3459 41010 4259 41040
rect 4609 41030 4639 41060
rect 4719 41030 4749 41060
rect 4829 41030 4859 41060
rect 4939 41030 4969 41060
rect 5049 41030 5079 41060
rect 5159 41030 5189 41060
rect 5269 41030 5299 41060
rect 5379 41030 5409 41060
rect 2509 40970 2539 41000
rect 2619 40970 2649 41000
rect 2729 40970 2759 41000
rect 2839 40970 2869 41000
rect 2949 40970 2979 41000
rect 3459 40990 3519 41010
rect 4609 41000 5409 41030
rect 2509 40940 3039 40970
rect 2979 40900 2989 40940
rect 3029 40900 3039 40940
rect 3459 40950 3469 40990
rect 3509 40950 3519 40990
rect 3459 40930 3519 40950
rect 5349 40980 5409 41000
rect 5349 40940 5359 40980
rect 5399 40940 5409 40980
rect 6019 40950 6049 40980
rect 6249 40950 6279 40980
rect 6359 40950 6389 40980
rect 6589 40950 6619 40980
rect 6699 40950 6729 40980
rect 6809 40950 6839 40980
rect 6919 40950 6949 40980
rect 7149 40950 7179 40980
rect 7259 40950 7289 40980
rect 7369 40950 7399 40980
rect 7479 40950 7509 40980
rect 7589 40950 7619 40980
rect 7699 40950 7729 40980
rect 7809 40950 7839 40980
rect 7919 40950 7949 40980
rect 8209 40950 8239 40980
rect 8319 40950 8349 40980
rect 8429 40950 8459 40980
rect 8539 40950 8569 40980
rect 8649 40950 8679 40980
rect 8759 40950 8789 40980
rect 8869 40950 8899 40980
rect 8979 40950 9009 40980
rect 9089 40950 9119 40980
rect 9199 40950 9229 40980
rect 9309 40950 9339 40980
rect 9419 40950 9449 40980
rect 9529 40950 9559 40980
rect 9639 40950 9669 40980
rect 9749 40950 9779 40980
rect 9859 40950 9889 40980
rect 5349 40920 5409 40940
rect 2979 40880 3039 40900
rect 2989 40660 3079 40680
rect 2989 40620 2999 40660
rect 3039 40620 3079 40660
rect 2989 40600 3079 40620
rect 2719 40560 2749 40590
rect 3049 40560 3079 40600
rect 3329 40530 3359 40560
rect 3439 40530 3469 40560
rect 3549 40530 3579 40560
rect 3659 40530 3689 40560
rect 3769 40530 3799 40560
rect 3879 40530 3909 40560
rect 3989 40530 4019 40560
rect 4099 40530 4129 40560
rect 4609 40530 4639 40560
rect 4719 40530 4749 40560
rect 4829 40530 4859 40560
rect 4939 40530 4969 40560
rect 5049 40530 5079 40560
rect 5159 40530 5189 40560
rect 5269 40530 5299 40560
rect 5379 40530 5409 40560
rect 6419 40520 6449 40550
rect 6529 40520 6559 40550
rect 6639 40520 6669 40550
rect 6749 40520 6779 40550
rect 6859 40520 6889 40550
rect 6969 40520 6999 40550
rect 7079 40520 7109 40550
rect 7189 40520 7219 40550
rect 7299 40520 7329 40550
rect 7409 40520 7439 40550
rect 7519 40520 7549 40550
rect 7629 40520 7659 40550
rect 7739 40520 7769 40550
rect 7849 40520 7879 40550
rect 7959 40520 7989 40550
rect 8069 40520 8099 40550
rect 8179 40520 8209 40550
rect 8289 40520 8319 40550
rect 8399 40520 8429 40550
rect 8509 40520 8539 40550
rect 8619 40520 8649 40550
rect 8729 40520 8759 40550
rect 8839 40520 8869 40550
rect 8949 40520 8979 40550
rect 9059 40520 9089 40550
rect 9169 40520 9199 40550
rect 9279 40520 9309 40550
rect 9389 40520 9419 40550
rect 9499 40520 9529 40550
rect 9609 40520 9639 40550
rect 9719 40520 9749 40550
rect 9829 40520 9859 40550
rect 6419 39980 6449 40020
rect 6349 39960 6449 39980
rect 6349 39920 6369 39960
rect 6409 39940 6449 39960
rect 6529 39940 6559 40020
rect 6639 39940 6669 40020
rect 6749 39940 6779 40020
rect 6859 39940 6889 40020
rect 6969 39940 6999 40020
rect 7079 39940 7109 40020
rect 7189 39940 7219 40020
rect 7299 39940 7329 40020
rect 7409 39940 7439 40020
rect 7519 39940 7549 40020
rect 7629 39940 7659 40020
rect 7739 39940 7769 40020
rect 7849 39940 7879 40020
rect 7959 39940 7989 40020
rect 8069 39940 8099 40020
rect 8179 39940 8209 40020
rect 8289 39940 8319 40020
rect 8399 39940 8429 40020
rect 8509 39940 8539 40020
rect 8619 39940 8649 40020
rect 8729 39940 8759 40020
rect 8839 39940 8869 40020
rect 8949 39940 8979 40020
rect 9059 39940 9089 40020
rect 9169 39940 9199 40020
rect 9279 39940 9309 40020
rect 9389 39940 9419 40020
rect 9499 39940 9529 40020
rect 9609 39940 9639 40020
rect 9719 39940 9749 40020
rect 9829 39940 9859 40020
rect 6409 39920 9859 39940
rect 6349 39900 9859 39920
rect 6419 39860 6449 39900
rect 6529 39860 6559 39900
rect 6639 39860 6669 39900
rect 6749 39860 6779 39900
rect 6859 39860 6889 39900
rect 6969 39860 6999 39900
rect 7079 39860 7109 39900
rect 7189 39860 7219 39900
rect 7299 39860 7329 39900
rect 7409 39860 7439 39900
rect 7519 39860 7549 39900
rect 7629 39860 7659 39900
rect 7739 39860 7769 39900
rect 7849 39860 7879 39900
rect 7959 39860 7989 39900
rect 8069 39860 8099 39900
rect 8179 39860 8209 39900
rect 8289 39860 8319 39900
rect 8399 39860 8429 39900
rect 8509 39860 8539 39900
rect 8619 39860 8649 39900
rect 8729 39860 8759 39900
rect 8839 39860 8869 39900
rect 8949 39860 8979 39900
rect 9059 39860 9089 39900
rect 9169 39860 9199 39900
rect 9279 39860 9309 39900
rect 9389 39860 9419 39900
rect 9499 39860 9529 39900
rect 9609 39860 9639 39900
rect 9719 39860 9749 39900
rect 9829 39860 9859 39900
rect 2719 39710 2749 39760
rect 3049 39730 3079 39760
rect 3329 39750 3359 39780
rect 3439 39750 3469 39780
rect 3549 39750 3579 39780
rect 3659 39750 3689 39780
rect 3769 39750 3799 39780
rect 3879 39750 3909 39780
rect 3989 39750 4019 39780
rect 4099 39750 4129 39780
rect 3329 39720 4129 39750
rect 4609 39750 4639 39780
rect 4719 39750 4749 39780
rect 4829 39750 4859 39780
rect 4939 39750 4969 39780
rect 5049 39750 5079 39780
rect 5159 39750 5189 39780
rect 5269 39750 5299 39780
rect 5379 39750 5409 39780
rect 4609 39720 5409 39750
rect 2719 39690 2809 39710
rect 2719 39650 2759 39690
rect 2799 39650 2809 39690
rect 2719 39630 2809 39650
rect 3329 39700 3389 39720
rect 3329 39660 3339 39700
rect 3379 39660 3389 39700
rect 3329 39640 3389 39660
rect 5349 39700 5409 39720
rect 5349 39660 5359 39700
rect 5399 39660 5409 39700
rect 5349 39640 5409 39660
rect 6419 39630 6449 39660
rect 6529 39630 6559 39660
rect 6639 39630 6669 39660
rect 6749 39630 6779 39660
rect 6859 39630 6889 39660
rect 6969 39630 6999 39660
rect 7079 39630 7109 39660
rect 7189 39630 7219 39660
rect 7299 39630 7329 39660
rect 7409 39630 7439 39660
rect 7519 39630 7549 39660
rect 7629 39630 7659 39660
rect 7739 39630 7769 39660
rect 7849 39630 7879 39660
rect 7959 39630 7989 39660
rect 8069 39630 8099 39660
rect 8179 39630 8209 39660
rect 8289 39630 8319 39660
rect 8399 39630 8429 39660
rect 8509 39630 8539 39660
rect 8619 39630 8649 39660
rect 8729 39630 8759 39660
rect 8839 39630 8869 39660
rect 8949 39630 8979 39660
rect 9059 39630 9089 39660
rect 9169 39630 9199 39660
rect 9279 39630 9309 39660
rect 9389 39630 9419 39660
rect 9499 39630 9529 39660
rect 9609 39630 9639 39660
rect 9719 39630 9749 39660
rect 9829 39630 9859 39660
rect 3840 37050 3870 37080
rect 3950 37050 3980 37080
rect 4060 37050 4090 37080
rect 4170 37050 4200 37080
rect 4280 37050 4310 37080
rect 4390 37050 4420 37080
rect 4650 37050 4680 37080
rect 4760 37050 4790 37080
rect 4870 37050 4900 37080
rect 4980 37050 5010 37080
rect 5090 37050 5120 37080
rect 5200 37050 5230 37080
rect 5530 37050 5560 37080
rect 5640 37050 5670 37080
rect 5750 37050 5780 37080
rect 5860 37050 5890 37080
rect 5970 37050 6000 37080
rect 6080 37050 6110 37080
rect 3840 35010 3870 36250
rect 3730 34990 3870 35010
rect 3950 34990 3980 36250
rect 4060 34990 4090 36250
rect 4170 34990 4200 36250
rect 4280 34990 4310 36250
rect 4390 34990 4420 36250
rect 4650 35010 4680 36250
rect 3730 34940 3760 34990
rect 3810 34940 4420 34990
rect 3730 34920 3870 34940
rect 3840 34690 3870 34920
rect 3950 34690 3980 34940
rect 4060 34690 4090 34940
rect 4170 34690 4200 34940
rect 4280 34690 4310 34940
rect 4390 34690 4420 34940
rect 4530 35000 4680 35010
rect 4530 34930 4560 35000
rect 4620 34990 4680 35000
rect 4760 34990 4790 36250
rect 4870 34990 4900 36250
rect 4980 34990 5010 36250
rect 5090 34990 5120 36250
rect 5200 34990 5230 36250
rect 4620 34940 5230 34990
rect 4620 34930 4680 34940
rect 4530 34920 4680 34930
rect 4650 34690 4680 34920
rect 4760 34690 4790 34940
rect 4870 34690 4900 34940
rect 4980 34690 5010 34940
rect 5090 34690 5120 34940
rect 5200 34690 5230 34940
rect 5530 34890 5560 36650
rect 5390 34870 5560 34890
rect 5640 34870 5670 36650
rect 5750 34870 5780 36650
rect 5860 34870 5890 36650
rect 5970 34870 6000 36650
rect 6080 34870 6110 36650
rect 6410 36590 6440 36620
rect 6520 36590 6550 36620
rect 6770 36590 6800 36620
rect 6880 36590 6910 36620
rect 7030 36590 7060 36620
rect 7140 36590 7170 36620
rect 7370 36590 7400 36620
rect 7480 36590 7510 36620
rect 7750 36590 7780 36620
rect 7860 36590 7890 36620
rect 8130 36590 8160 36620
rect 8240 36590 8270 36620
rect 8510 36590 8540 36620
rect 8620 36590 8650 36620
rect 8850 36590 8880 36620
rect 8960 36590 8990 36620
rect 9110 36590 9140 36620
rect 9220 36590 9250 36620
rect 9450 36590 9480 36620
rect 9560 36590 9590 36620
rect 9830 36590 9860 36620
rect 9940 36590 9970 36620
rect 10210 36590 10240 36620
rect 10320 36590 10350 36620
rect 10590 36590 10620 36620
rect 10700 36590 10730 36620
rect 5390 34820 5420 34870
rect 5470 34820 6110 34870
rect 6410 34860 6440 36390
rect 5390 34800 5560 34820
rect 5530 34760 5560 34800
rect 5640 34760 5670 34820
rect 5750 34760 5780 34820
rect 5860 34760 5890 34820
rect 5970 34760 6000 34820
rect 6080 34760 6110 34820
rect 6320 34850 6440 34860
rect 6520 34850 6550 36390
rect 7370 36370 7400 36390
rect 7480 36370 7510 36390
rect 7370 36340 7510 36370
rect 6770 34870 6800 36190
rect 6320 34810 6340 34850
rect 6380 34810 6550 34850
rect 6320 34800 6440 34810
rect 6410 34760 6440 34800
rect 6520 34760 6550 34810
rect 6710 34850 6800 34870
rect 6880 34850 6910 36190
rect 6710 34810 6720 34850
rect 6760 34820 6910 34850
rect 6760 34810 6800 34820
rect 6710 34790 6800 34810
rect 6770 34750 6800 34790
rect 6880 34750 6910 34820
rect 7030 34750 7060 36190
rect 7140 34750 7170 36190
rect 7370 34850 7400 36340
rect 7280 34840 7400 34850
rect 7280 34800 7300 34840
rect 7340 34800 7400 34840
rect 7280 34790 7400 34800
rect 7370 34750 7400 34790
rect 7480 34750 7510 36340
rect 7750 36370 7780 36390
rect 7860 36370 7890 36390
rect 7750 36340 7890 36370
rect 7750 34850 7780 36340
rect 7660 34840 7780 34850
rect 7660 34800 7680 34840
rect 7720 34800 7780 34840
rect 7660 34790 7780 34800
rect 7750 34750 7780 34790
rect 7860 34750 7890 36340
rect 8130 36370 8160 36390
rect 8240 36370 8270 36390
rect 8130 36340 8270 36370
rect 8130 34850 8160 36340
rect 8040 34840 8160 34850
rect 8040 34800 8060 34840
rect 8100 34800 8160 34840
rect 8040 34790 8160 34800
rect 8130 34750 8160 34790
rect 8240 34750 8270 36340
rect 8510 36370 8540 36390
rect 8620 36370 8650 36390
rect 8510 36340 8650 36370
rect 8510 34850 8540 36340
rect 8420 34840 8540 34850
rect 8420 34800 8440 34840
rect 8480 34800 8540 34840
rect 8420 34790 8540 34800
rect 8510 34750 8540 34790
rect 8620 34750 8650 36340
rect 9450 36370 9480 36390
rect 9560 36370 9590 36390
rect 9450 36340 9590 36370
rect 8850 34860 8880 36190
rect 8790 34840 8880 34860
rect 8960 34840 8990 36190
rect 9110 34970 9140 36190
rect 9050 34950 9140 34970
rect 9050 34910 9060 34950
rect 9100 34940 9140 34950
rect 9220 34940 9250 36190
rect 9100 34910 9250 34940
rect 9050 34890 9140 34910
rect 8790 34800 8800 34840
rect 8840 34810 8990 34840
rect 8840 34800 8880 34810
rect 8790 34780 8880 34800
rect 8850 34750 8880 34780
rect 8960 34750 8990 34810
rect 9110 34750 9140 34890
rect 9220 34750 9250 34910
rect 9450 34850 9480 36340
rect 9360 34840 9480 34850
rect 9360 34800 9380 34840
rect 9420 34800 9480 34840
rect 9360 34790 9480 34800
rect 9450 34750 9480 34790
rect 9560 34750 9590 36340
rect 9830 36370 9860 36390
rect 9940 36370 9970 36390
rect 9830 36340 9970 36370
rect 9830 34850 9860 36340
rect 9740 34840 9860 34850
rect 9740 34800 9760 34840
rect 9800 34800 9860 34840
rect 9740 34790 9860 34800
rect 9830 34750 9860 34790
rect 9940 34750 9970 36340
rect 10210 36370 10240 36390
rect 10320 36370 10350 36390
rect 10210 36340 10350 36370
rect 10210 34850 10240 36340
rect 10120 34840 10240 34850
rect 10120 34800 10140 34840
rect 10180 34800 10240 34840
rect 10120 34790 10240 34800
rect 10210 34750 10240 34790
rect 10320 34750 10350 36340
rect 10590 36370 10620 36390
rect 10700 36370 10730 36390
rect 10590 36340 10730 36370
rect 10590 34850 10620 36340
rect 10500 34840 10620 34850
rect 10500 34800 10520 34840
rect 10560 34800 10620 34840
rect 10500 34790 10620 34800
rect 10590 34750 10620 34790
rect 10700 34750 10730 36340
rect 15410 36110 15520 36120
rect 15410 36070 15460 36110
rect 15500 36070 15520 36110
rect 17530 36080 17560 36110
rect 17780 36080 17810 36110
rect 18100 36080 18130 36110
rect 18470 36080 18500 36110
rect 18720 36080 18750 36110
rect 19040 36080 19070 36110
rect 19830 36100 19860 36130
rect 20080 36100 20110 36130
rect 15410 36060 15520 36070
rect 15410 35970 15440 36060
rect 15520 35970 15550 36000
rect 16530 35840 16560 35870
rect 16640 35840 16670 35870
rect 16750 35840 16780 35870
rect 16860 35840 16890 35870
rect 16970 35840 17000 35870
rect 17080 35840 17110 35870
rect 15410 35740 15440 35770
rect 15520 35640 15550 35770
rect 15520 35630 15660 35640
rect 15520 35570 15570 35630
rect 15640 35570 15660 35630
rect 15520 35560 15660 35570
rect 16530 35510 16560 35610
rect 16430 35500 16560 35510
rect 16640 35500 16670 35610
rect 16750 35500 16780 35610
rect 16860 35500 16890 35610
rect 16970 35500 17000 35610
rect 17080 35500 17110 35610
rect 19370 36010 19400 36040
rect 16430 35490 17110 35500
rect 16430 35430 16450 35490
rect 16510 35440 17110 35490
rect 17530 35500 17560 35580
rect 17780 35500 17810 35580
rect 18100 35500 18130 35580
rect 17530 35490 17640 35500
rect 17530 35450 17580 35490
rect 17620 35450 17640 35490
rect 17530 35440 17640 35450
rect 17700 35490 17810 35500
rect 17700 35450 17720 35490
rect 17760 35450 17810 35490
rect 17700 35440 17810 35450
rect 18020 35490 18130 35500
rect 18020 35450 18040 35490
rect 18080 35450 18130 35490
rect 18020 35440 18130 35450
rect 18470 35500 18500 35580
rect 18720 35500 18750 35580
rect 19040 35500 19070 35580
rect 18470 35490 18580 35500
rect 18470 35450 18520 35490
rect 18560 35450 18580 35490
rect 18470 35440 18580 35450
rect 18640 35490 18750 35500
rect 18640 35450 18660 35490
rect 18700 35450 18750 35490
rect 18640 35440 18750 35450
rect 18960 35490 19070 35500
rect 18960 35450 18980 35490
rect 19020 35450 19070 35490
rect 18960 35440 19070 35450
rect 16510 35430 16560 35440
rect 16430 35410 16560 35430
rect 16530 35350 16560 35410
rect 16640 35350 16670 35440
rect 16750 35350 16780 35440
rect 16860 35350 16890 35440
rect 16970 35350 17000 35440
rect 17080 35350 17110 35440
rect 6410 34230 6440 34260
rect 6520 34230 6550 34260
rect 17820 35200 17930 35210
rect 17420 35160 17450 35190
rect 17820 35160 17870 35200
rect 17910 35160 17930 35200
rect 18360 35160 18390 35190
rect 18760 35160 18790 35190
rect 17820 35150 17930 35160
rect 17820 35110 17850 35150
rect 17420 34910 17450 34960
rect 22490 36080 22520 36110
rect 22740 36080 22770 36110
rect 23060 36080 23090 36110
rect 23430 36080 23460 36110
rect 23680 36080 23710 36110
rect 24000 36080 24030 36110
rect 24790 36100 24820 36130
rect 25040 36100 25070 36130
rect 21100 36010 21130 36040
rect 19830 35500 19860 35600
rect 20080 35530 20110 35600
rect 19750 35490 19860 35500
rect 19750 35450 19770 35490
rect 19810 35450 19860 35490
rect 20000 35520 20110 35530
rect 20000 35480 20020 35520
rect 20060 35480 20110 35520
rect 20000 35470 20110 35480
rect 19750 35440 19860 35450
rect 19830 35150 19860 35180
rect 20080 35150 20110 35180
rect 19370 34970 19400 35010
rect 18360 34910 18390 34960
rect 18760 34910 18790 34960
rect 17420 34900 17530 34910
rect 17420 34860 17470 34900
rect 17510 34860 17530 34900
rect 17820 34880 17850 34910
rect 18360 34900 18470 34910
rect 17420 34850 17530 34860
rect 18360 34860 18410 34900
rect 18450 34860 18470 34900
rect 18360 34850 18470 34860
rect 18680 34900 18790 34910
rect 18680 34860 18700 34900
rect 18740 34860 18790 34900
rect 19310 34950 19400 34970
rect 21490 35840 21520 35870
rect 21600 35840 21630 35870
rect 21710 35840 21740 35870
rect 21820 35840 21850 35870
rect 21930 35840 21960 35870
rect 22040 35840 22070 35870
rect 21490 35500 21520 35610
rect 21600 35500 21630 35610
rect 21710 35500 21740 35610
rect 21820 35500 21850 35610
rect 21930 35500 21960 35610
rect 22040 35500 22070 35610
rect 24330 36010 24360 36040
rect 21410 35490 22070 35500
rect 21410 35450 21430 35490
rect 21470 35450 22070 35490
rect 21410 35440 22070 35450
rect 22490 35500 22520 35580
rect 22740 35500 22770 35580
rect 23060 35500 23090 35580
rect 22490 35490 22600 35500
rect 22490 35450 22540 35490
rect 22580 35450 22600 35490
rect 22490 35440 22600 35450
rect 22660 35490 22770 35500
rect 22660 35450 22680 35490
rect 22720 35450 22770 35490
rect 22660 35440 22770 35450
rect 22980 35490 23090 35500
rect 22980 35450 23000 35490
rect 23040 35450 23090 35490
rect 22980 35440 23090 35450
rect 23430 35500 23460 35580
rect 23680 35500 23710 35580
rect 24000 35500 24030 35580
rect 23430 35490 23540 35500
rect 23430 35450 23480 35490
rect 23520 35450 23540 35490
rect 23430 35440 23540 35450
rect 23600 35490 23710 35500
rect 23600 35450 23620 35490
rect 23660 35450 23710 35490
rect 23600 35440 23710 35450
rect 23920 35490 24030 35500
rect 23920 35450 23940 35490
rect 23980 35450 24030 35490
rect 23920 35440 24030 35450
rect 21490 35350 21520 35440
rect 21600 35350 21630 35440
rect 21710 35350 21740 35440
rect 21820 35350 21850 35440
rect 21930 35350 21960 35440
rect 22040 35350 22070 35440
rect 20900 34960 21000 34980
rect 19310 34910 19320 34950
rect 19360 34910 19400 34950
rect 19310 34890 19400 34910
rect 18680 34850 18790 34860
rect 19370 34850 19400 34890
rect 17640 34640 17670 34670
rect 18100 34640 18130 34670
rect 18580 34640 18610 34670
rect 19040 34640 19070 34670
rect 16530 34420 16560 34450
rect 16640 34420 16670 34450
rect 16750 34420 16780 34450
rect 16860 34420 16890 34450
rect 16970 34420 17000 34450
rect 17080 34420 17110 34450
rect 19830 34830 19860 34950
rect 19730 34810 19860 34830
rect 20080 34820 20110 34950
rect 20900 34900 20920 34960
rect 20980 34950 21000 34960
rect 21100 34950 21130 35010
rect 20980 34910 21130 34950
rect 20980 34900 21000 34910
rect 20900 34880 21000 34900
rect 21100 34850 21130 34910
rect 19730 34750 19750 34810
rect 19810 34750 19860 34810
rect 20000 34810 20110 34820
rect 20000 34770 20020 34810
rect 20060 34770 20110 34810
rect 20000 34760 20110 34770
rect 19730 34730 19860 34750
rect 19750 34660 19860 34670
rect 19750 34620 19770 34660
rect 19810 34620 19860 34660
rect 19750 34610 19860 34620
rect 19830 34570 19860 34610
rect 17640 34370 17670 34440
rect 18100 34370 18130 34440
rect 17640 34360 17750 34370
rect 17640 34320 17690 34360
rect 17730 34320 17750 34360
rect 17640 34310 17750 34320
rect 18020 34360 18130 34370
rect 18020 34320 18040 34360
rect 18080 34320 18130 34360
rect 18020 34310 18130 34320
rect 18580 34370 18610 34440
rect 19040 34370 19070 34440
rect 19370 34420 19400 34450
rect 22780 35200 22890 35210
rect 22380 35160 22410 35190
rect 22780 35160 22830 35200
rect 22870 35160 22890 35200
rect 23320 35160 23350 35190
rect 23720 35160 23750 35190
rect 22780 35150 22890 35160
rect 22780 35110 22810 35150
rect 22380 34910 22410 34960
rect 24790 35500 24820 35600
rect 25040 35530 25070 35600
rect 24710 35490 24820 35500
rect 24710 35450 24730 35490
rect 24770 35450 24820 35490
rect 24960 35520 25070 35530
rect 24960 35480 24980 35520
rect 25020 35480 25070 35520
rect 24960 35470 25070 35480
rect 24710 35440 24820 35450
rect 24790 35150 24820 35180
rect 25040 35150 25070 35180
rect 24330 34970 24360 35010
rect 23320 34910 23350 34960
rect 23720 34910 23750 34960
rect 22380 34900 22490 34910
rect 22380 34860 22430 34900
rect 22470 34860 22490 34900
rect 22780 34880 22810 34910
rect 23320 34900 23430 34910
rect 22380 34850 22490 34860
rect 23320 34860 23370 34900
rect 23410 34860 23430 34900
rect 23320 34850 23430 34860
rect 23640 34900 23750 34910
rect 23640 34860 23660 34900
rect 23700 34860 23750 34900
rect 24270 34950 24360 34970
rect 24270 34910 24280 34950
rect 24320 34910 24360 34950
rect 24270 34890 24360 34910
rect 23640 34850 23750 34860
rect 24330 34850 24360 34890
rect 22600 34640 22630 34670
rect 23060 34640 23090 34670
rect 23540 34640 23570 34670
rect 24000 34640 24030 34670
rect 21100 34420 21130 34450
rect 21490 34420 21520 34450
rect 21600 34420 21630 34450
rect 21710 34420 21740 34450
rect 21820 34420 21850 34450
rect 21930 34420 21960 34450
rect 22040 34420 22070 34450
rect 24790 34830 24820 34950
rect 24690 34810 24820 34830
rect 25040 34820 25070 34950
rect 24690 34750 24710 34810
rect 24770 34750 24820 34810
rect 24960 34810 25070 34820
rect 24960 34770 24980 34810
rect 25020 34770 25070 34810
rect 24960 34760 25070 34770
rect 24690 34730 24820 34750
rect 24710 34660 24820 34670
rect 24710 34620 24730 34660
rect 24770 34620 24820 34660
rect 24710 34610 24820 34620
rect 24790 34570 24820 34610
rect 22600 34370 22630 34440
rect 23060 34370 23090 34440
rect 18580 34360 18690 34370
rect 18580 34320 18630 34360
rect 18670 34320 18690 34360
rect 18580 34310 18690 34320
rect 18960 34360 19070 34370
rect 18960 34320 18980 34360
rect 19020 34320 19070 34360
rect 19830 34340 19860 34370
rect 22600 34360 22710 34370
rect 18960 34310 19070 34320
rect 22600 34320 22650 34360
rect 22690 34320 22710 34360
rect 22600 34310 22710 34320
rect 22980 34360 23090 34370
rect 22980 34320 23000 34360
rect 23040 34320 23090 34360
rect 22980 34310 23090 34320
rect 23540 34370 23570 34440
rect 24000 34370 24030 34440
rect 24330 34420 24360 34450
rect 23540 34360 23650 34370
rect 23540 34320 23590 34360
rect 23630 34320 23650 34360
rect 23540 34310 23650 34320
rect 23920 34360 24030 34370
rect 23920 34320 23940 34360
rect 23980 34320 24030 34360
rect 24790 34340 24820 34370
rect 23920 34310 24030 34320
rect 6770 34220 6800 34250
rect 6880 34220 6910 34250
rect 7030 34170 7060 34250
rect 7140 34210 7170 34250
rect 7370 34220 7400 34250
rect 7480 34220 7510 34250
rect 7750 34220 7780 34250
rect 7860 34220 7890 34250
rect 8130 34220 8160 34250
rect 8240 34220 8270 34250
rect 8510 34220 8540 34250
rect 8620 34220 8650 34250
rect 8850 34220 8880 34250
rect 8960 34220 8990 34250
rect 9110 34220 9140 34250
rect 9220 34220 9250 34250
rect 9450 34220 9480 34250
rect 9560 34220 9590 34250
rect 9830 34220 9860 34250
rect 9940 34220 9970 34250
rect 10210 34220 10240 34250
rect 10320 34220 10350 34250
rect 10590 34220 10620 34250
rect 10700 34220 10730 34250
rect 7140 34190 7230 34210
rect 7140 34170 7180 34190
rect 7030 34150 7180 34170
rect 7220 34150 7230 34190
rect 7030 34140 7230 34150
rect 7030 34110 7060 34140
rect 7140 34130 7230 34140
rect 7140 34110 7170 34130
rect 5530 33730 5560 33760
rect 5640 33730 5670 33760
rect 5750 33730 5780 33760
rect 5860 33730 5890 33760
rect 5970 33730 6000 33760
rect 6080 33730 6110 33760
rect 3840 33660 3870 33690
rect 3950 33660 3980 33690
rect 4060 33660 4090 33690
rect 4170 33660 4200 33690
rect 4280 33660 4310 33690
rect 4390 33660 4420 33690
rect 4650 33660 4680 33690
rect 4760 33660 4790 33690
rect 4870 33660 4900 33690
rect 4980 33660 5010 33690
rect 5090 33660 5120 33690
rect 5200 33660 5230 33690
rect 14068 32380 14178 32390
rect 14068 32340 14118 32380
rect 14158 32340 14178 32380
rect 14068 32330 14178 32340
rect 13958 32240 13988 32270
rect 14068 32240 14098 32330
rect 14178 32240 14208 32270
rect 13958 31950 13988 32040
rect 14068 32010 14098 32040
rect 13958 31940 14068 31950
rect 13958 31900 14008 31940
rect 14048 31900 14068 31940
rect 13958 31890 14068 31900
rect 14178 31900 14208 32040
rect 17530 32020 17560 32050
rect 17780 32020 17810 32050
rect 18100 32020 18130 32050
rect 18470 32020 18500 32050
rect 18720 32020 18750 32050
rect 19040 32020 19070 32050
rect 20090 32020 20120 32050
rect 20340 32020 20370 32050
rect 14178 31890 14288 31900
rect 14178 31850 14228 31890
rect 14268 31850 14288 31890
rect 14178 31840 14288 31850
rect 16530 31780 16560 31810
rect 16640 31780 16670 31810
rect 16750 31780 16780 31810
rect 16860 31780 16890 31810
rect 16970 31780 17000 31810
rect 17080 31780 17110 31810
rect 14178 31660 14208 31690
rect 2240 31600 2270 31630
rect 2350 31600 2380 31630
rect 2460 31600 2490 31630
rect 2570 31600 2600 31630
rect 2680 31600 2710 31630
rect 2790 31600 2820 31630
rect 3050 31600 3080 31630
rect 3160 31600 3190 31630
rect 3270 31600 3300 31630
rect 3380 31600 3410 31630
rect 3490 31600 3520 31630
rect 3600 31600 3630 31630
rect 3930 31600 3960 31630
rect 4040 31600 4070 31630
rect 4150 31600 4180 31630
rect 4260 31600 4290 31630
rect 4370 31600 4400 31630
rect 4480 31600 4510 31630
rect 4790 31600 4820 31630
rect 4900 31600 4930 31630
rect 5010 31600 5040 31630
rect 5120 31600 5150 31630
rect 5230 31600 5260 31630
rect 5340 31600 5370 31630
rect 5650 31600 5680 31630
rect 5760 31600 5790 31630
rect 5870 31600 5900 31630
rect 5980 31600 6010 31630
rect 6090 31600 6120 31630
rect 6200 31600 6230 31630
rect 16530 31470 16560 31550
rect 16430 31450 16560 31470
rect 16430 31390 16450 31450
rect 16510 31440 16560 31450
rect 16640 31440 16670 31550
rect 16750 31440 16780 31550
rect 16860 31440 16890 31550
rect 16970 31440 17000 31550
rect 17080 31440 17110 31550
rect 19370 31950 19400 31980
rect 19630 31950 19660 31980
rect 16510 31390 17110 31440
rect 16430 31380 17110 31390
rect 17530 31440 17560 31520
rect 17780 31440 17810 31520
rect 18100 31440 18130 31520
rect 17530 31430 17640 31440
rect 17530 31390 17580 31430
rect 17620 31390 17640 31430
rect 17530 31380 17640 31390
rect 17700 31430 17810 31440
rect 17700 31390 17720 31430
rect 17760 31390 17810 31430
rect 17700 31380 17810 31390
rect 18020 31430 18130 31440
rect 18020 31390 18040 31430
rect 18080 31390 18130 31430
rect 18020 31380 18130 31390
rect 18470 31440 18500 31520
rect 18720 31440 18750 31520
rect 19040 31440 19070 31520
rect 18470 31430 18580 31440
rect 18470 31390 18520 31430
rect 18560 31390 18580 31430
rect 18470 31380 18580 31390
rect 18640 31430 18750 31440
rect 18640 31390 18660 31430
rect 18700 31390 18750 31430
rect 18640 31380 18750 31390
rect 18960 31430 19070 31440
rect 18960 31390 18980 31430
rect 19020 31390 19070 31430
rect 18960 31380 19070 31390
rect 16430 31370 16560 31380
rect 14178 31320 14208 31360
rect 14098 31310 14208 31320
rect 14098 31270 14118 31310
rect 14158 31270 14208 31310
rect 16530 31290 16560 31370
rect 16640 31290 16670 31380
rect 16750 31290 16780 31380
rect 16860 31290 16890 31380
rect 16970 31290 17000 31380
rect 17080 31290 17110 31380
rect 6470 31240 6500 31270
rect 6580 31240 6610 31270
rect 6830 31240 6860 31270
rect 6940 31240 6970 31270
rect 7090 31240 7120 31270
rect 7200 31240 7230 31270
rect 7430 31240 7460 31270
rect 7540 31240 7570 31270
rect 7810 31240 7840 31270
rect 7920 31240 7950 31270
rect 8190 31240 8220 31270
rect 8300 31240 8330 31270
rect 8570 31240 8600 31270
rect 8680 31240 8710 31270
rect 8910 31240 8940 31270
rect 9020 31240 9050 31270
rect 9170 31240 9200 31270
rect 9280 31240 9310 31270
rect 9510 31240 9540 31270
rect 9620 31240 9650 31270
rect 9890 31240 9920 31270
rect 10000 31240 10030 31270
rect 10270 31240 10300 31270
rect 10380 31240 10410 31270
rect 10650 31240 10680 31270
rect 10760 31240 10790 31270
rect 11030 31240 11060 31270
rect 11140 31240 11170 31270
rect 14098 31260 14208 31270
rect 2240 30760 2270 30800
rect 2350 30760 2380 30800
rect 2460 30760 2490 30800
rect 2570 30760 2600 30800
rect 2680 30760 2710 30800
rect 2790 30760 2820 30800
rect 3050 30760 3080 30800
rect 3160 30760 3190 30800
rect 3270 30760 3300 30800
rect 3380 30760 3410 30800
rect 3490 30760 3520 30800
rect 3600 30760 3630 30800
rect 2130 30740 2820 30760
rect 2130 30690 2160 30740
rect 2210 30690 2820 30740
rect 2130 30670 2820 30690
rect 2930 30740 3630 30760
rect 2930 30680 2960 30740
rect 3020 30680 3630 30740
rect 2930 30670 3630 30680
rect 2240 30440 2270 30670
rect 2350 30440 2380 30670
rect 2460 30440 2490 30670
rect 2570 30440 2600 30670
rect 2680 30440 2710 30670
rect 2790 30440 2820 30670
rect 3050 30440 3080 30670
rect 3160 30440 3190 30670
rect 3270 30440 3300 30670
rect 3380 30440 3410 30670
rect 3490 30440 3520 30670
rect 3600 30440 3630 30670
rect 3930 30610 3960 31200
rect 4040 30610 4070 31200
rect 4150 30610 4180 31200
rect 4260 30610 4290 31200
rect 4370 30610 4400 31200
rect 4480 30610 4510 31200
rect 4790 30620 4820 31200
rect 3790 30600 4510 30610
rect 3790 30560 3820 30600
rect 3860 30560 4510 30600
rect 3790 30550 4510 30560
rect 4660 30610 4820 30620
rect 4900 30610 4930 31200
rect 5010 30610 5040 31200
rect 5120 30610 5150 31200
rect 5230 30610 5260 31200
rect 5340 30610 5370 31200
rect 5650 30620 5680 31200
rect 4660 30560 4680 30610
rect 4730 30560 5370 30610
rect 4660 30550 5370 30560
rect 5520 30610 5680 30620
rect 5760 30610 5790 31200
rect 5870 30610 5900 31200
rect 5980 30610 6010 31200
rect 6090 30610 6120 31200
rect 6200 30610 6230 31200
rect 6470 31020 6500 31040
rect 6580 31020 6610 31040
rect 6470 30990 6610 31020
rect 6470 30710 6500 30990
rect 6380 30700 6500 30710
rect 6380 30660 6400 30700
rect 6440 30660 6500 30700
rect 6380 30650 6500 30660
rect 6470 30610 6500 30650
rect 6580 30610 6610 30990
rect 7430 31020 7460 31040
rect 7540 31020 7570 31040
rect 7430 30990 7570 31020
rect 6830 30720 6860 30840
rect 6770 30700 6860 30720
rect 6770 30660 6780 30700
rect 6820 30690 6860 30700
rect 6940 30690 6970 30840
rect 6820 30660 6970 30690
rect 6770 30640 6860 30660
rect 5520 30560 5540 30610
rect 5590 30560 6230 30610
rect 5520 30550 6230 30560
rect 3930 30510 3960 30550
rect 4040 30510 4070 30550
rect 4150 30510 4180 30550
rect 4260 30510 4290 30550
rect 4370 30510 4400 30550
rect 4480 30510 4510 30550
rect 4790 30510 4820 30550
rect 4900 30510 4930 30550
rect 5010 30510 5040 30550
rect 5120 30510 5150 30550
rect 5230 30510 5260 30550
rect 5340 30510 5370 30550
rect 5650 30510 5680 30550
rect 5760 30510 5790 30550
rect 5870 30510 5900 30550
rect 5980 30510 6010 30550
rect 6090 30510 6120 30550
rect 6200 30510 6230 30550
rect 6830 30600 6860 30640
rect 6940 30600 6970 30660
rect 7090 30600 7120 30840
rect 7200 30600 7230 30840
rect 7430 30700 7460 30990
rect 7540 30700 7570 30990
rect 7810 31020 7840 31040
rect 7920 31020 7950 31040
rect 7810 30990 7950 31020
rect 7810 30700 7840 30990
rect 7340 30690 7460 30700
rect 7340 30650 7360 30690
rect 7400 30650 7460 30690
rect 7340 30640 7460 30650
rect 7720 30690 7840 30700
rect 7720 30650 7740 30690
rect 7780 30650 7840 30690
rect 7720 30640 7840 30650
rect 7430 30600 7460 30640
rect 7540 30600 7570 30640
rect 7810 30600 7840 30640
rect 7920 30600 7950 30990
rect 8190 31020 8220 31040
rect 8300 31020 8330 31040
rect 8190 30990 8330 31020
rect 8190 30700 8220 30990
rect 8100 30690 8220 30700
rect 8100 30650 8120 30690
rect 8160 30650 8220 30690
rect 8100 30640 8220 30650
rect 8190 30600 8220 30640
rect 8300 30600 8330 30990
rect 8570 31020 8600 31040
rect 8680 31020 8710 31040
rect 8570 30990 8710 31020
rect 8570 30700 8600 30990
rect 8480 30690 8600 30700
rect 8480 30650 8500 30690
rect 8540 30650 8600 30690
rect 8480 30640 8600 30650
rect 8570 30600 8600 30640
rect 8680 30600 8710 30990
rect 9510 31020 9540 31040
rect 9620 31020 9650 31040
rect 9510 30990 9650 31020
rect 8910 30710 8940 30840
rect 8850 30690 8940 30710
rect 9020 30690 9050 30840
rect 9170 30820 9200 30840
rect 9110 30800 9200 30820
rect 9110 30760 9120 30800
rect 9160 30790 9200 30800
rect 9280 30790 9310 30840
rect 9160 30760 9310 30790
rect 9110 30740 9200 30760
rect 8850 30650 8860 30690
rect 8900 30660 9050 30690
rect 8900 30650 8940 30660
rect 8850 30630 8940 30650
rect 8910 30600 8940 30630
rect 9020 30600 9050 30660
rect 9170 30600 9200 30740
rect 9280 30600 9310 30760
rect 9510 30700 9540 30990
rect 9420 30690 9540 30700
rect 9420 30650 9440 30690
rect 9480 30650 9540 30690
rect 9420 30640 9540 30650
rect 9510 30600 9540 30640
rect 9620 30600 9650 30990
rect 9890 31020 9920 31040
rect 10000 31020 10030 31040
rect 9890 30990 10030 31020
rect 9890 30700 9920 30990
rect 9800 30690 9920 30700
rect 9800 30650 9820 30690
rect 9860 30650 9920 30690
rect 9800 30640 9920 30650
rect 9890 30600 9920 30640
rect 10000 30600 10030 30990
rect 10270 31020 10300 31040
rect 10380 31020 10410 31040
rect 10270 30990 10410 31020
rect 10270 30700 10300 30990
rect 10180 30690 10300 30700
rect 10180 30650 10200 30690
rect 10240 30650 10300 30690
rect 10180 30640 10300 30650
rect 10270 30600 10300 30640
rect 10380 30600 10410 30990
rect 10650 31020 10680 31040
rect 10760 31020 10790 31040
rect 10650 30990 10790 31020
rect 10650 30700 10680 30990
rect 10560 30690 10680 30700
rect 10560 30650 10580 30690
rect 10620 30650 10680 30690
rect 10560 30640 10680 30650
rect 10650 30600 10680 30640
rect 10760 30600 10790 30990
rect 11030 31020 11060 31040
rect 11140 31020 11170 31040
rect 11030 30990 11170 31020
rect 11030 30700 11060 30990
rect 10940 30690 11060 30700
rect 10940 30650 10960 30690
rect 11000 30650 11060 30690
rect 10940 30640 11060 30650
rect 11030 30600 11060 30640
rect 11140 30600 11170 30990
rect 6470 30080 6500 30110
rect 6580 30080 6610 30110
rect 17820 31140 17930 31150
rect 17420 31100 17450 31130
rect 17820 31100 17870 31140
rect 17910 31100 17930 31140
rect 18360 31100 18390 31130
rect 18760 31100 18790 31130
rect 17820 31090 17930 31100
rect 17820 31050 17850 31090
rect 17420 30850 17450 30900
rect 22550 32010 22580 32040
rect 22800 32010 22830 32040
rect 23120 32010 23150 32040
rect 23490 32010 23520 32040
rect 23740 32010 23770 32040
rect 24060 32010 24090 32040
rect 25050 32030 25080 32060
rect 25300 32030 25330 32060
rect 21160 31950 21190 31980
rect 20090 31440 20120 31520
rect 20340 31450 20370 31520
rect 20010 31430 20120 31440
rect 20010 31390 20030 31430
rect 20070 31390 20120 31430
rect 20260 31440 20370 31450
rect 20260 31400 20280 31440
rect 20320 31400 20370 31440
rect 20260 31390 20370 31400
rect 20010 31380 20120 31390
rect 20090 31090 20120 31120
rect 20340 31090 20370 31120
rect 19370 30910 19400 30950
rect 19630 30910 19660 30950
rect 18360 30850 18390 30900
rect 18760 30850 18790 30900
rect 17420 30840 17530 30850
rect 17420 30800 17470 30840
rect 17510 30800 17530 30840
rect 17820 30820 17850 30850
rect 18360 30840 18470 30850
rect 17420 30790 17530 30800
rect 18360 30800 18410 30840
rect 18450 30800 18470 30840
rect 18360 30790 18470 30800
rect 18680 30840 18790 30850
rect 18680 30800 18700 30840
rect 18740 30800 18790 30840
rect 19310 30890 19400 30910
rect 19310 30850 19320 30890
rect 19360 30850 19400 30890
rect 19310 30830 19400 30850
rect 19570 30890 19660 30910
rect 21550 31770 21580 31800
rect 21660 31770 21690 31800
rect 21770 31770 21800 31800
rect 21880 31770 21910 31800
rect 21990 31770 22020 31800
rect 22100 31770 22130 31800
rect 21550 31430 21580 31540
rect 21660 31430 21690 31540
rect 21770 31430 21800 31540
rect 21880 31430 21910 31540
rect 21990 31430 22020 31540
rect 22100 31430 22130 31540
rect 24390 31940 24420 31970
rect 24650 31940 24680 31970
rect 21470 31420 22130 31430
rect 21470 31380 21490 31420
rect 21530 31380 22130 31420
rect 21470 31370 22130 31380
rect 22550 31430 22580 31510
rect 22800 31430 22830 31510
rect 23120 31430 23150 31510
rect 22550 31420 22660 31430
rect 22550 31380 22600 31420
rect 22640 31380 22660 31420
rect 22550 31370 22660 31380
rect 22720 31420 22830 31430
rect 22720 31380 22740 31420
rect 22780 31380 22830 31420
rect 22720 31370 22830 31380
rect 23040 31420 23150 31430
rect 23040 31380 23060 31420
rect 23100 31380 23150 31420
rect 23040 31370 23150 31380
rect 23490 31430 23520 31510
rect 23740 31430 23770 31510
rect 24060 31430 24090 31510
rect 23490 31420 23600 31430
rect 23490 31380 23540 31420
rect 23580 31380 23600 31420
rect 23490 31370 23600 31380
rect 23660 31420 23770 31430
rect 23660 31380 23680 31420
rect 23720 31380 23770 31420
rect 23660 31370 23770 31380
rect 23980 31420 24090 31430
rect 23980 31380 24000 31420
rect 24040 31380 24090 31420
rect 23980 31370 24090 31380
rect 21550 31280 21580 31370
rect 21660 31280 21690 31370
rect 21770 31280 21800 31370
rect 21880 31280 21910 31370
rect 21990 31280 22020 31370
rect 22100 31280 22130 31370
rect 20960 30900 21060 30920
rect 19570 30850 19580 30890
rect 19620 30850 19660 30890
rect 19570 30830 19660 30850
rect 18680 30790 18790 30800
rect 19370 30790 19400 30830
rect 19630 30790 19660 30830
rect 17640 30580 17670 30610
rect 18100 30580 18130 30610
rect 18580 30580 18610 30610
rect 19040 30580 19070 30610
rect 16530 30360 16560 30390
rect 16640 30360 16670 30390
rect 16750 30360 16780 30390
rect 16860 30360 16890 30390
rect 16970 30360 17000 30390
rect 17080 30360 17110 30390
rect 20090 30770 20120 30890
rect 19990 30750 20120 30770
rect 20340 30760 20370 30890
rect 20960 30840 20980 30900
rect 21040 30890 21060 30900
rect 21160 30890 21190 30950
rect 21040 30850 21190 30890
rect 21040 30840 21060 30850
rect 20960 30820 21060 30840
rect 21160 30790 21190 30850
rect 19990 30690 20010 30750
rect 20070 30690 20120 30750
rect 20260 30750 20370 30760
rect 20260 30710 20280 30750
rect 20320 30710 20370 30750
rect 20260 30700 20370 30710
rect 19990 30670 20120 30690
rect 20010 30600 20120 30610
rect 20010 30560 20030 30600
rect 20070 30560 20120 30600
rect 20010 30550 20120 30560
rect 20090 30510 20120 30550
rect 17640 30310 17670 30380
rect 18100 30310 18130 30380
rect 17640 30300 17750 30310
rect 17640 30260 17690 30300
rect 17730 30260 17750 30300
rect 17640 30250 17750 30260
rect 18020 30300 18130 30310
rect 18020 30260 18040 30300
rect 18080 30260 18130 30300
rect 18020 30250 18130 30260
rect 18580 30310 18610 30380
rect 19040 30310 19070 30380
rect 19370 30360 19400 30390
rect 19630 30360 19660 30390
rect 21160 30360 21190 30390
rect 22840 31130 22950 31140
rect 22440 31090 22470 31120
rect 22840 31090 22890 31130
rect 22930 31090 22950 31130
rect 23380 31090 23410 31120
rect 23780 31090 23810 31120
rect 22840 31080 22950 31090
rect 22840 31040 22870 31080
rect 22440 30840 22470 30890
rect 25050 31430 25080 31530
rect 25300 31460 25330 31530
rect 24970 31420 25080 31430
rect 24970 31380 24990 31420
rect 25030 31380 25080 31420
rect 25220 31450 25330 31460
rect 25220 31410 25240 31450
rect 25280 31410 25330 31450
rect 25220 31400 25330 31410
rect 24970 31370 25080 31380
rect 25050 31080 25080 31110
rect 25300 31080 25330 31110
rect 24390 30900 24420 30940
rect 24650 30900 24680 30940
rect 23380 30840 23410 30890
rect 23780 30840 23810 30890
rect 22440 30830 22550 30840
rect 22440 30790 22490 30830
rect 22530 30790 22550 30830
rect 22840 30810 22870 30840
rect 23380 30830 23490 30840
rect 22440 30780 22550 30790
rect 23380 30790 23430 30830
rect 23470 30790 23490 30830
rect 23380 30780 23490 30790
rect 23700 30830 23810 30840
rect 23700 30790 23720 30830
rect 23760 30790 23810 30830
rect 24330 30880 24420 30900
rect 24330 30840 24340 30880
rect 24380 30840 24420 30880
rect 24330 30820 24420 30840
rect 24590 30880 24680 30900
rect 24590 30840 24600 30880
rect 24640 30840 24680 30880
rect 24590 30820 24680 30840
rect 23700 30780 23810 30790
rect 24390 30780 24420 30820
rect 24650 30780 24680 30820
rect 22660 30570 22690 30600
rect 23120 30570 23150 30600
rect 23600 30570 23630 30600
rect 24060 30570 24090 30600
rect 21550 30350 21580 30380
rect 21660 30350 21690 30380
rect 21770 30350 21800 30380
rect 21880 30350 21910 30380
rect 21990 30350 22020 30380
rect 22100 30350 22130 30380
rect 25050 30760 25080 30880
rect 24950 30740 25080 30760
rect 25300 30750 25330 30880
rect 24950 30680 24970 30740
rect 25030 30680 25080 30740
rect 25220 30740 25330 30750
rect 25220 30700 25240 30740
rect 25280 30700 25330 30740
rect 25220 30690 25330 30700
rect 24950 30660 25080 30680
rect 24970 30590 25080 30600
rect 24970 30550 24990 30590
rect 25030 30550 25080 30590
rect 24970 30540 25080 30550
rect 25050 30500 25080 30540
rect 18580 30300 18690 30310
rect 18580 30260 18630 30300
rect 18670 30260 18690 30300
rect 18580 30250 18690 30260
rect 18960 30300 19070 30310
rect 18960 30260 18980 30300
rect 19020 30260 19070 30300
rect 20090 30280 20120 30310
rect 22660 30300 22690 30370
rect 23120 30300 23150 30370
rect 22660 30290 22770 30300
rect 18960 30250 19070 30260
rect 22660 30250 22710 30290
rect 22750 30250 22770 30290
rect 22660 30240 22770 30250
rect 23040 30290 23150 30300
rect 23040 30250 23060 30290
rect 23100 30250 23150 30290
rect 23040 30240 23150 30250
rect 23600 30300 23630 30370
rect 24060 30300 24090 30370
rect 24390 30350 24420 30380
rect 24650 30350 24680 30380
rect 23600 30290 23710 30300
rect 23600 30250 23650 30290
rect 23690 30250 23710 30290
rect 23600 30240 23710 30250
rect 23980 30290 24090 30300
rect 23980 30250 24000 30290
rect 24040 30250 24090 30290
rect 25050 30270 25080 30300
rect 23980 30240 24090 30250
rect 6830 30070 6860 30100
rect 6940 30070 6970 30100
rect 7090 30020 7120 30100
rect 7200 30060 7230 30100
rect 7430 30070 7460 30100
rect 7540 30070 7570 30100
rect 7810 30070 7840 30100
rect 7920 30070 7950 30100
rect 8190 30070 8220 30100
rect 8300 30070 8330 30100
rect 8570 30070 8600 30100
rect 8680 30070 8710 30100
rect 8910 30070 8940 30100
rect 9020 30070 9050 30100
rect 9170 30070 9200 30100
rect 9280 30070 9310 30100
rect 9510 30070 9540 30100
rect 9620 30070 9650 30100
rect 9890 30070 9920 30100
rect 10000 30070 10030 30100
rect 10270 30070 10300 30100
rect 10380 30070 10410 30100
rect 10650 30070 10680 30100
rect 10760 30070 10790 30100
rect 11030 30070 11060 30100
rect 11140 30070 11170 30100
rect 7200 30040 7290 30060
rect 7200 30020 7240 30040
rect 7090 30000 7240 30020
rect 7280 30000 7290 30040
rect 7090 29990 7290 30000
rect 7090 29960 7120 29990
rect 7200 29980 7290 29990
rect 7200 29960 7230 29980
rect 3930 29480 3960 29510
rect 4040 29480 4070 29510
rect 4150 29480 4180 29510
rect 4260 29480 4290 29510
rect 4370 29480 4400 29510
rect 4480 29480 4510 29510
rect 4790 29480 4820 29510
rect 4900 29480 4930 29510
rect 5010 29480 5040 29510
rect 5120 29480 5150 29510
rect 5230 29480 5260 29510
rect 5340 29480 5370 29510
rect 5650 29480 5680 29510
rect 5760 29480 5790 29510
rect 5870 29480 5900 29510
rect 5980 29480 6010 29510
rect 6090 29480 6120 29510
rect 6200 29480 6230 29510
rect 2240 29410 2270 29440
rect 2350 29410 2380 29440
rect 2460 29410 2490 29440
rect 2570 29410 2600 29440
rect 2680 29410 2710 29440
rect 2790 29410 2820 29440
rect 3050 29410 3080 29440
rect 3160 29410 3190 29440
rect 3270 29410 3300 29440
rect 3380 29410 3410 29440
rect 3490 29410 3520 29440
rect 3600 29410 3630 29440
rect 7390 26490 7420 26520
rect 7500 26490 7530 26520
rect 7920 26490 7950 26520
rect 8030 26490 8060 26520
rect 8550 26500 8580 26530
rect 8700 26500 8730 26530
rect 8930 26500 8960 26530
rect 9290 26500 9320 26530
rect 9400 26500 9430 26530
rect 9630 26500 9660 26530
rect 9740 26500 9770 26530
rect 9890 26500 9920 26530
rect 10000 26500 10030 26530
rect 10230 26500 10260 26530
rect 10340 26500 10370 26530
rect 10620 26500 10650 26530
rect 10730 26500 10760 26530
rect 10880 26500 10910 26530
rect 10990 26500 11020 26530
rect 11220 26500 11250 26530
rect 11330 26500 11360 26530
rect 11620 26500 11650 26530
rect 11730 26500 11760 26530
rect 11880 26500 11910 26530
rect 11990 26500 12020 26530
rect 12220 26500 12250 26530
rect 12330 26500 12360 26530
rect 12600 26500 12630 26530
rect 12710 26500 12740 26530
rect 12950 26500 12980 26530
rect 13180 26500 13210 26530
rect 13290 26500 13320 26530
rect 13520 26500 13550 26530
rect 13630 26500 13660 26530
rect 13740 26500 13770 26530
rect 13850 26500 13880 26530
rect 14080 26500 14110 26530
rect 14190 26500 14220 26530
rect 14300 26500 14330 26530
rect 14410 26500 14440 26530
rect 14520 26500 14550 26530
rect 14630 26500 14660 26530
rect 14740 26500 14770 26530
rect 14850 26500 14880 26530
rect 15140 26500 15170 26530
rect 15250 26500 15280 26530
rect 15360 26500 15390 26530
rect 15470 26500 15500 26530
rect 15580 26500 15610 26530
rect 15690 26500 15720 26530
rect 15800 26500 15830 26530
rect 15910 26500 15940 26530
rect 16020 26500 16050 26530
rect 16130 26500 16160 26530
rect 16240 26500 16270 26530
rect 16350 26500 16380 26530
rect 16460 26500 16490 26530
rect 16570 26500 16600 26530
rect 16680 26500 16710 26530
rect 16790 26500 16820 26530
rect 17090 26500 17120 26530
rect 17200 26500 17230 26530
rect 17310 26500 17340 26530
rect 17420 26500 17450 26530
rect 17530 26500 17560 26530
rect 17640 26500 17670 26530
rect 17750 26500 17780 26530
rect 17860 26500 17890 26530
rect 17970 26500 18000 26530
rect 18080 26500 18110 26530
rect 18190 26500 18220 26530
rect 18300 26500 18330 26530
rect 18410 26500 18440 26530
rect 18520 26500 18550 26530
rect 18630 26500 18660 26530
rect 18740 26500 18770 26530
rect 18850 26500 18880 26530
rect 18960 26500 18990 26530
rect 19070 26500 19100 26530
rect 19180 26500 19210 26530
rect 19290 26500 19320 26530
rect 19400 26500 19430 26530
rect 19510 26500 19540 26530
rect 19620 26500 19650 26530
rect 19730 26500 19760 26530
rect 19840 26500 19870 26530
rect 19950 26500 19980 26530
rect 20060 26500 20090 26530
rect 20170 26500 20200 26530
rect 20280 26500 20310 26530
rect 20390 26500 20420 26530
rect 20500 26500 20530 26530
rect 7390 25210 7420 25990
rect 7270 25190 7420 25210
rect 7270 25130 7290 25190
rect 7350 25130 7420 25190
rect 7270 25110 7420 25130
rect 7390 24620 7420 25110
rect 7500 24620 7530 25990
rect 7920 25580 7950 25990
rect 7800 25560 7950 25580
rect 7800 25500 7820 25560
rect 7880 25500 7950 25560
rect 7800 25480 7950 25500
rect 7390 24590 7530 24620
rect 7390 24570 7420 24590
rect 7500 24570 7530 24590
rect 7920 24620 7950 25480
rect 8030 24620 8060 25990
rect 8550 24960 8580 26000
rect 8480 24940 8580 24960
rect 8480 24900 8500 24940
rect 8540 24900 8580 24940
rect 8480 24880 8580 24900
rect 8700 24880 8730 26000
rect 8930 24960 8960 26000
rect 9290 24960 9320 26000
rect 8860 24940 8960 24960
rect 8860 24900 8880 24940
rect 8920 24900 8960 24940
rect 9200 24950 9320 24960
rect 9200 24910 9220 24950
rect 9260 24910 9320 24950
rect 9200 24900 9320 24910
rect 8860 24880 8960 24900
rect 8550 24760 8580 24880
rect 8630 24860 8730 24880
rect 8630 24820 8650 24860
rect 8690 24820 8730 24860
rect 8930 24830 8960 24880
rect 8630 24800 8730 24820
rect 8700 24760 8730 24800
rect 7920 24590 8060 24620
rect 7920 24570 7950 24590
rect 8030 24570 8060 24590
rect 7390 24340 7420 24370
rect 7500 24340 7530 24370
rect 7920 24340 7950 24370
rect 8030 24340 8060 24370
rect 8930 24600 8960 24630
rect 9290 24560 9320 24900
rect 9400 24560 9430 26000
rect 9630 25960 9660 26000
rect 9740 25960 9770 26000
rect 9630 25950 9770 25960
rect 9630 25910 9680 25950
rect 9720 25910 9770 25950
rect 9630 25900 9770 25910
rect 9890 25960 9920 26000
rect 10000 25960 10030 26000
rect 9890 25950 10030 25960
rect 9890 25910 9940 25950
rect 9980 25910 10030 25950
rect 9890 25900 10030 25910
rect 9630 25060 9770 25070
rect 9630 25020 9680 25060
rect 9720 25020 9770 25060
rect 9630 25010 9770 25020
rect 9630 24960 9660 25010
rect 9570 24940 9660 24960
rect 9740 24940 9770 25010
rect 9570 24900 9580 24940
rect 9620 24910 9770 24940
rect 9620 24900 9660 24910
rect 9570 24880 9660 24900
rect 9630 24760 9660 24880
rect 9740 24760 9770 24910
rect 9890 25060 10030 25070
rect 9890 25020 9940 25060
rect 9980 25020 10030 25060
rect 9890 25010 10030 25020
rect 9890 24860 9920 25010
rect 9830 24840 9920 24860
rect 9830 24800 9840 24840
rect 9880 24800 9920 24840
rect 9830 24780 9920 24800
rect 9890 24760 9920 24780
rect 10000 24760 10030 25010
rect 10230 24960 10260 26000
rect 10140 24950 10260 24960
rect 10140 24910 10160 24950
rect 10200 24910 10260 24950
rect 10140 24900 10260 24910
rect 10230 24800 10260 24900
rect 10340 24800 10370 26000
rect 10620 25960 10650 26000
rect 10730 25960 10760 26000
rect 10620 25950 10760 25960
rect 10620 25910 10670 25950
rect 10710 25910 10760 25950
rect 10620 25900 10760 25910
rect 10880 25960 10910 26000
rect 10990 25960 11020 26000
rect 10880 25950 11020 25960
rect 10880 25910 10930 25950
rect 10970 25910 11020 25950
rect 10880 25900 11020 25910
rect 10620 25060 10760 25070
rect 10620 25020 10670 25060
rect 10710 25020 10760 25060
rect 10620 25010 10760 25020
rect 10620 24960 10650 25010
rect 10560 24940 10650 24960
rect 10730 24940 10760 25010
rect 10560 24900 10570 24940
rect 10610 24910 10760 24940
rect 10610 24900 10650 24910
rect 10560 24880 10650 24900
rect 10230 24760 10370 24800
rect 10620 24760 10650 24880
rect 10730 24760 10760 24910
rect 10880 25060 11020 25070
rect 10880 25020 10930 25060
rect 10970 25020 11020 25060
rect 10880 25010 11020 25020
rect 10880 24860 10910 25010
rect 10820 24840 10910 24860
rect 10990 24840 11020 25010
rect 11220 24960 11250 26000
rect 11130 24950 11250 24960
rect 11130 24910 11150 24950
rect 11190 24910 11250 24950
rect 11130 24900 11250 24910
rect 10820 24800 10830 24840
rect 10870 24810 11020 24840
rect 10870 24800 10910 24810
rect 10820 24780 10910 24800
rect 10880 24760 10910 24780
rect 10990 24760 11020 24810
rect 11220 24800 11250 24900
rect 11330 24800 11360 26000
rect 11620 25960 11650 26000
rect 11730 25960 11760 26000
rect 11620 25950 11760 25960
rect 11620 25910 11670 25950
rect 11710 25910 11760 25950
rect 11620 25900 11760 25910
rect 11880 25960 11910 26000
rect 11990 25960 12020 26000
rect 11880 25950 12020 25960
rect 11880 25910 11930 25950
rect 11970 25910 12020 25950
rect 11880 25900 12020 25910
rect 11620 25060 11760 25070
rect 11620 25020 11670 25060
rect 11710 25020 11760 25060
rect 11620 25010 11760 25020
rect 11620 24960 11650 25010
rect 11560 24940 11650 24960
rect 11560 24900 11570 24940
rect 11610 24900 11650 24940
rect 11560 24880 11650 24900
rect 11220 24770 11360 24800
rect 10230 24560 10260 24760
rect 10340 24560 10370 24760
rect 11220 24560 11250 24770
rect 11330 24560 11360 24770
rect 11620 24760 11650 24880
rect 11730 24760 11760 25010
rect 11880 25060 12020 25070
rect 11880 25020 11930 25060
rect 11970 25020 12020 25060
rect 11880 25010 12020 25020
rect 11880 24860 11910 25010
rect 11820 24840 11910 24860
rect 11820 24800 11830 24840
rect 11870 24800 11910 24840
rect 11820 24780 11910 24800
rect 11880 24760 11910 24780
rect 11990 24760 12020 25010
rect 12220 24960 12250 26000
rect 12130 24950 12250 24960
rect 12130 24910 12150 24950
rect 12190 24910 12250 24950
rect 12130 24900 12250 24910
rect 12220 24780 12250 24900
rect 12330 24780 12360 26000
rect 12600 24960 12630 26000
rect 12510 24950 12630 24960
rect 12510 24910 12530 24950
rect 12570 24910 12630 24950
rect 12510 24900 12630 24910
rect 12220 24750 12360 24780
rect 12220 24560 12250 24750
rect 12330 24560 12360 24750
rect 12600 24780 12630 24900
rect 12710 24780 12740 26000
rect 12950 24960 12980 26000
rect 13180 25940 13210 26000
rect 13290 25940 13320 26000
rect 13180 25930 13320 25940
rect 13180 25890 13230 25930
rect 13270 25890 13320 25930
rect 13180 25880 13320 25890
rect 13520 25940 13550 26000
rect 13630 25940 13660 26000
rect 13520 25930 13660 25940
rect 13520 25890 13570 25930
rect 13610 25890 13660 25930
rect 13520 25880 13660 25890
rect 13740 25940 13770 26000
rect 13850 25940 13880 26000
rect 13740 25930 13880 25940
rect 13740 25890 13790 25930
rect 13830 25890 13880 25930
rect 14080 25960 14110 26000
rect 14190 25960 14220 26000
rect 14080 25950 14220 25960
rect 14080 25910 14130 25950
rect 14170 25910 14220 25950
rect 14080 25900 14220 25910
rect 14300 25960 14330 26000
rect 14410 25960 14440 26000
rect 14300 25950 14440 25960
rect 14300 25910 14350 25950
rect 14390 25910 14440 25950
rect 14300 25900 14440 25910
rect 14520 25960 14550 26000
rect 14630 25960 14660 26000
rect 14520 25950 14660 25960
rect 14520 25910 14570 25950
rect 14610 25910 14660 25950
rect 14520 25900 14660 25910
rect 14740 25960 14770 26000
rect 14850 25960 14880 26000
rect 14740 25950 14880 25960
rect 14740 25910 14790 25950
rect 14830 25910 14880 25950
rect 14740 25900 14880 25910
rect 15140 25960 15170 26000
rect 15250 25960 15280 26000
rect 15140 25950 15280 25960
rect 15140 25910 15190 25950
rect 15230 25910 15280 25950
rect 15140 25900 15280 25910
rect 15360 25960 15390 26000
rect 15470 25960 15500 26000
rect 15360 25950 15500 25960
rect 15360 25910 15410 25950
rect 15450 25910 15500 25950
rect 15360 25900 15500 25910
rect 15580 25960 15610 26000
rect 15690 25960 15720 26000
rect 15580 25950 15720 25960
rect 15580 25910 15630 25950
rect 15670 25910 15720 25950
rect 15580 25900 15720 25910
rect 15800 25960 15830 26000
rect 15910 25960 15940 26000
rect 15800 25950 15940 25960
rect 15800 25910 15850 25950
rect 15890 25910 15940 25950
rect 15800 25900 15940 25910
rect 16020 25960 16050 26000
rect 16130 25960 16160 26000
rect 16020 25950 16160 25960
rect 16020 25910 16070 25950
rect 16110 25910 16160 25950
rect 16020 25900 16160 25910
rect 16240 25960 16270 26000
rect 16350 25960 16380 26000
rect 16240 25950 16380 25960
rect 16240 25910 16290 25950
rect 16330 25910 16380 25950
rect 16240 25900 16380 25910
rect 16460 25960 16490 26000
rect 16570 25960 16600 26000
rect 16460 25950 16600 25960
rect 16460 25910 16510 25950
rect 16550 25910 16600 25950
rect 16460 25900 16600 25910
rect 16680 25960 16710 26000
rect 16790 25960 16820 26000
rect 16680 25950 16820 25960
rect 16680 25910 16730 25950
rect 16770 25910 16820 25950
rect 16680 25900 16820 25910
rect 17090 25960 17120 26000
rect 17200 25960 17230 26000
rect 17090 25950 17230 25960
rect 17090 25910 17140 25950
rect 17180 25910 17230 25950
rect 17090 25900 17230 25910
rect 17310 25960 17340 26000
rect 17420 25960 17450 26000
rect 17310 25950 17450 25960
rect 17310 25910 17360 25950
rect 17400 25910 17450 25950
rect 17310 25900 17450 25910
rect 17530 25960 17560 26000
rect 17640 25960 17670 26000
rect 17530 25950 17670 25960
rect 17530 25910 17580 25950
rect 17620 25910 17670 25950
rect 17530 25900 17670 25910
rect 17750 25960 17780 26000
rect 17860 25960 17890 26000
rect 17750 25950 17890 25960
rect 17750 25910 17800 25950
rect 17840 25910 17890 25950
rect 17750 25900 17890 25910
rect 17970 25960 18000 26000
rect 18080 25960 18110 26000
rect 17970 25950 18110 25960
rect 17970 25910 18020 25950
rect 18060 25910 18110 25950
rect 17970 25900 18110 25910
rect 18190 25960 18220 26000
rect 18300 25960 18330 26000
rect 18190 25950 18330 25960
rect 18190 25910 18240 25950
rect 18280 25910 18330 25950
rect 18190 25900 18330 25910
rect 18410 25960 18440 26000
rect 18520 25960 18550 26000
rect 18410 25950 18550 25960
rect 18410 25910 18460 25950
rect 18500 25910 18550 25950
rect 18410 25900 18550 25910
rect 18630 25960 18660 26000
rect 18740 25960 18770 26000
rect 18630 25950 18770 25960
rect 18630 25910 18680 25950
rect 18720 25910 18770 25950
rect 18630 25900 18770 25910
rect 18850 25960 18880 26000
rect 18960 25960 18990 26000
rect 18850 25950 18990 25960
rect 18850 25910 18900 25950
rect 18940 25910 18990 25950
rect 18850 25900 18990 25910
rect 19070 25960 19100 26000
rect 19180 25960 19210 26000
rect 19070 25950 19210 25960
rect 19070 25910 19120 25950
rect 19160 25910 19210 25950
rect 19070 25900 19210 25910
rect 19290 25960 19320 26000
rect 19400 25960 19430 26000
rect 19290 25950 19430 25960
rect 19290 25910 19340 25950
rect 19380 25910 19430 25950
rect 19290 25900 19430 25910
rect 19510 25960 19540 26000
rect 19620 25960 19650 26000
rect 19510 25950 19650 25960
rect 19510 25910 19560 25950
rect 19600 25910 19650 25950
rect 19510 25900 19650 25910
rect 19730 25960 19760 26000
rect 19840 25960 19870 26000
rect 19730 25950 19870 25960
rect 19730 25910 19780 25950
rect 19820 25910 19870 25950
rect 19730 25900 19870 25910
rect 19950 25960 19980 26000
rect 20060 25960 20090 26000
rect 19950 25950 20090 25960
rect 19950 25910 20000 25950
rect 20040 25910 20090 25950
rect 19950 25900 20090 25910
rect 20170 25960 20200 26000
rect 20280 25960 20310 26000
rect 20170 25950 20310 25960
rect 20170 25910 20220 25950
rect 20260 25910 20310 25950
rect 20170 25900 20310 25910
rect 20390 25960 20420 26000
rect 20500 25960 20530 26000
rect 20390 25950 20530 25960
rect 20390 25910 20440 25950
rect 20480 25910 20530 25950
rect 20390 25900 20530 25910
rect 13740 25880 13880 25890
rect 14080 25060 14220 25070
rect 13180 25040 13320 25050
rect 13180 25000 13230 25040
rect 13270 25000 13320 25040
rect 13180 24990 13320 25000
rect 13180 24960 13210 24990
rect 12890 24940 12980 24960
rect 12890 24900 12900 24940
rect 12940 24900 12980 24940
rect 12890 24880 12980 24900
rect 13120 24940 13210 24960
rect 13120 24900 13130 24940
rect 13170 24920 13210 24940
rect 13290 24920 13320 24990
rect 13520 25040 13660 25050
rect 13520 25000 13570 25040
rect 13610 25000 13660 25040
rect 13520 24990 13660 25000
rect 13520 24960 13550 24990
rect 13170 24900 13320 24920
rect 13120 24880 13320 24900
rect 13460 24940 13550 24960
rect 13460 24900 13470 24940
rect 13510 24920 13550 24940
rect 13630 24920 13660 24990
rect 13740 25040 13880 25050
rect 13740 25000 13790 25040
rect 13830 25000 13880 25040
rect 13740 24990 13880 25000
rect 13740 24920 13770 24990
rect 13850 24920 13880 24990
rect 14080 25020 14130 25060
rect 14170 25020 14220 25060
rect 14080 25010 14220 25020
rect 14080 24960 14110 25010
rect 13510 24900 13880 24920
rect 13460 24880 13880 24900
rect 14020 24940 14110 24960
rect 14020 24900 14030 24940
rect 14070 24920 14110 24940
rect 14190 24920 14220 25010
rect 14300 25060 14440 25070
rect 14300 25020 14350 25060
rect 14390 25020 14440 25060
rect 14300 25010 14440 25020
rect 14300 24920 14330 25010
rect 14410 24920 14440 25010
rect 14520 25060 14660 25070
rect 14520 25020 14570 25060
rect 14610 25020 14660 25060
rect 14520 25010 14660 25020
rect 14520 24920 14550 25010
rect 14630 24920 14660 25010
rect 14740 25060 14880 25070
rect 14740 25020 14790 25060
rect 14830 25020 14880 25060
rect 14740 25010 14880 25020
rect 14740 24920 14770 25010
rect 14850 24920 14880 25010
rect 15140 25060 15280 25070
rect 15140 25020 15190 25060
rect 15230 25020 15280 25060
rect 15140 25010 15280 25020
rect 15140 24960 15170 25010
rect 14070 24900 14880 24920
rect 14020 24880 14880 24900
rect 15080 24940 15170 24960
rect 15080 24900 15090 24940
rect 15130 24920 15170 24940
rect 15250 24920 15280 25010
rect 15360 25060 15500 25070
rect 15360 25020 15410 25060
rect 15450 25020 15500 25060
rect 15360 25010 15500 25020
rect 15360 24920 15390 25010
rect 15470 24920 15500 25010
rect 15580 25060 15720 25070
rect 15580 25020 15630 25060
rect 15670 25020 15720 25060
rect 15580 25010 15720 25020
rect 15580 24920 15610 25010
rect 15690 24920 15720 25010
rect 15800 25060 15940 25070
rect 15800 25020 15850 25060
rect 15890 25020 15940 25060
rect 15800 25010 15940 25020
rect 15800 24920 15830 25010
rect 15910 24920 15940 25010
rect 16020 25060 16160 25070
rect 16020 25020 16070 25060
rect 16110 25020 16160 25060
rect 16020 25010 16160 25020
rect 16020 24920 16050 25010
rect 16130 24920 16160 25010
rect 16240 25060 16380 25070
rect 16240 25020 16290 25060
rect 16330 25020 16380 25060
rect 16240 25010 16380 25020
rect 16240 24920 16270 25010
rect 16350 24920 16380 25010
rect 16460 25060 16600 25070
rect 16460 25020 16510 25060
rect 16550 25020 16600 25060
rect 16460 25010 16600 25020
rect 16460 24920 16490 25010
rect 16570 24920 16600 25010
rect 16680 25060 16820 25070
rect 16680 25020 16730 25060
rect 16770 25020 16820 25060
rect 16680 25010 16820 25020
rect 16680 24920 16710 25010
rect 16790 24920 16820 25010
rect 17090 25060 17230 25070
rect 17090 25020 17140 25060
rect 17180 25020 17230 25060
rect 17090 25010 17230 25020
rect 17090 24960 17120 25010
rect 15130 24900 16820 24920
rect 15080 24880 16820 24900
rect 17020 24940 17120 24960
rect 17020 24900 17040 24940
rect 17080 24920 17120 24940
rect 17200 24920 17230 25010
rect 17310 25060 17450 25070
rect 17310 25020 17360 25060
rect 17400 25020 17450 25060
rect 17310 25010 17450 25020
rect 17310 24920 17340 25010
rect 17420 24920 17450 25010
rect 17530 25060 17670 25070
rect 17530 25020 17580 25060
rect 17620 25020 17670 25060
rect 17530 25010 17670 25020
rect 17530 24920 17560 25010
rect 17640 24920 17670 25010
rect 17750 25060 17890 25070
rect 17750 25020 17800 25060
rect 17840 25020 17890 25060
rect 17750 25010 17890 25020
rect 17750 24920 17780 25010
rect 17860 24920 17890 25010
rect 17970 25060 18110 25070
rect 17970 25020 18020 25060
rect 18060 25020 18110 25060
rect 17970 25010 18110 25020
rect 17970 24920 18000 25010
rect 18080 24920 18110 25010
rect 18190 25060 18330 25070
rect 18190 25020 18240 25060
rect 18280 25020 18330 25060
rect 18190 25010 18330 25020
rect 18190 24920 18220 25010
rect 18300 24920 18330 25010
rect 18410 25060 18550 25070
rect 18410 25020 18460 25060
rect 18500 25020 18550 25060
rect 18410 25010 18550 25020
rect 18410 24920 18440 25010
rect 18520 24920 18550 25010
rect 18630 25060 18770 25070
rect 18630 25020 18680 25060
rect 18720 25020 18770 25060
rect 18630 25010 18770 25020
rect 18630 24920 18660 25010
rect 18740 24920 18770 25010
rect 18850 25060 18990 25070
rect 18850 25020 18900 25060
rect 18940 25020 18990 25060
rect 18850 25010 18990 25020
rect 18850 24920 18880 25010
rect 18960 24920 18990 25010
rect 19070 25060 19210 25070
rect 19070 25020 19120 25060
rect 19160 25020 19210 25060
rect 19070 25010 19210 25020
rect 19070 24920 19100 25010
rect 19180 24920 19210 25010
rect 19290 25060 19430 25070
rect 19290 25020 19340 25060
rect 19380 25020 19430 25060
rect 19290 25010 19430 25020
rect 19290 24920 19320 25010
rect 19400 24920 19430 25010
rect 19510 25060 19650 25070
rect 19510 25020 19560 25060
rect 19600 25020 19650 25060
rect 19510 25010 19650 25020
rect 19510 24920 19540 25010
rect 19620 24920 19650 25010
rect 19730 25060 19870 25070
rect 19730 25020 19780 25060
rect 19820 25020 19870 25060
rect 19730 25010 19870 25020
rect 19730 24920 19760 25010
rect 19840 24920 19870 25010
rect 19950 25060 20090 25070
rect 19950 25020 20000 25060
rect 20040 25020 20090 25060
rect 19950 25010 20090 25020
rect 19950 24920 19980 25010
rect 20060 24920 20090 25010
rect 20170 25060 20310 25070
rect 20170 25020 20220 25060
rect 20260 25020 20310 25060
rect 20170 25010 20310 25020
rect 20170 24920 20200 25010
rect 20280 24920 20310 25010
rect 20390 25060 20530 25070
rect 20390 25020 20440 25060
rect 20480 25020 20530 25060
rect 20390 25010 20530 25020
rect 20390 24920 20420 25010
rect 20500 24920 20530 25010
rect 17080 24900 20530 24920
rect 17020 24880 20530 24900
rect 12950 24840 12980 24880
rect 13180 24840 13210 24880
rect 13290 24840 13320 24880
rect 13520 24840 13550 24880
rect 13630 24840 13660 24880
rect 13740 24840 13770 24880
rect 13850 24840 13880 24880
rect 14080 24840 14110 24880
rect 14190 24840 14220 24880
rect 14300 24840 14330 24880
rect 14410 24840 14440 24880
rect 14520 24840 14550 24880
rect 14630 24840 14660 24880
rect 14740 24840 14770 24880
rect 14850 24840 14880 24880
rect 15140 24840 15170 24880
rect 15250 24840 15280 24880
rect 15360 24840 15390 24880
rect 15470 24840 15500 24880
rect 15580 24840 15610 24880
rect 15690 24840 15720 24880
rect 15800 24840 15830 24880
rect 15910 24840 15940 24880
rect 16020 24840 16050 24880
rect 16130 24840 16160 24880
rect 16240 24840 16270 24880
rect 16350 24840 16380 24880
rect 16460 24840 16490 24880
rect 16570 24840 16600 24880
rect 16680 24840 16710 24880
rect 16790 24840 16820 24880
rect 17090 24840 17120 24880
rect 17200 24840 17230 24880
rect 17310 24840 17340 24880
rect 17420 24840 17450 24880
rect 17530 24840 17560 24880
rect 17640 24840 17670 24880
rect 17750 24840 17780 24880
rect 17860 24840 17890 24880
rect 17970 24840 18000 24880
rect 18080 24840 18110 24880
rect 18190 24840 18220 24880
rect 18300 24840 18330 24880
rect 18410 24840 18440 24880
rect 18520 24840 18550 24880
rect 18630 24840 18660 24880
rect 18740 24840 18770 24880
rect 18850 24840 18880 24880
rect 18960 24840 18990 24880
rect 19070 24840 19100 24880
rect 19180 24840 19210 24880
rect 19290 24840 19320 24880
rect 19400 24840 19430 24880
rect 19510 24840 19540 24880
rect 19620 24840 19650 24880
rect 19730 24840 19760 24880
rect 19840 24840 19870 24880
rect 19950 24840 19980 24880
rect 20060 24840 20090 24880
rect 20170 24840 20200 24880
rect 20280 24840 20310 24880
rect 20390 24840 20420 24880
rect 20500 24840 20530 24880
rect 12600 24750 12740 24780
rect 12600 24560 12630 24750
rect 12710 24560 12740 24750
rect 12950 24610 12980 24640
rect 13180 24610 13210 24640
rect 13290 24610 13320 24640
rect 13520 24610 13550 24640
rect 13630 24610 13660 24640
rect 13740 24610 13770 24640
rect 13850 24610 13880 24640
rect 14080 24610 14110 24640
rect 14190 24610 14220 24640
rect 14300 24610 14330 24640
rect 14410 24610 14440 24640
rect 14520 24610 14550 24640
rect 14630 24610 14660 24640
rect 14740 24610 14770 24640
rect 14850 24610 14880 24640
rect 15140 24610 15170 24640
rect 15250 24610 15280 24640
rect 15360 24610 15390 24640
rect 15470 24610 15500 24640
rect 15580 24610 15610 24640
rect 15690 24610 15720 24640
rect 15800 24610 15830 24640
rect 15910 24610 15940 24640
rect 16020 24610 16050 24640
rect 16130 24610 16160 24640
rect 16240 24610 16270 24640
rect 16350 24610 16380 24640
rect 16460 24610 16490 24640
rect 16570 24610 16600 24640
rect 16680 24610 16710 24640
rect 16790 24610 16820 24640
rect 17090 24610 17120 24640
rect 17200 24610 17230 24640
rect 17310 24610 17340 24640
rect 17420 24610 17450 24640
rect 17530 24610 17560 24640
rect 17640 24610 17670 24640
rect 17750 24610 17780 24640
rect 17860 24610 17890 24640
rect 17970 24610 18000 24640
rect 18080 24610 18110 24640
rect 18190 24610 18220 24640
rect 18300 24610 18330 24640
rect 18410 24610 18440 24640
rect 18520 24610 18550 24640
rect 18630 24610 18660 24640
rect 18740 24610 18770 24640
rect 18850 24610 18880 24640
rect 18960 24610 18990 24640
rect 19070 24610 19100 24640
rect 19180 24610 19210 24640
rect 19290 24610 19320 24640
rect 19400 24610 19430 24640
rect 19510 24610 19540 24640
rect 19620 24610 19650 24640
rect 19730 24610 19760 24640
rect 19840 24610 19870 24640
rect 19950 24610 19980 24640
rect 20060 24610 20090 24640
rect 20170 24610 20200 24640
rect 20280 24610 20310 24640
rect 20390 24610 20420 24640
rect 20500 24610 20530 24640
rect 8550 24330 8580 24360
rect 8700 24330 8730 24360
rect 9290 24330 9320 24360
rect 9400 24330 9430 24360
rect 9630 24330 9660 24360
rect 9740 24330 9770 24360
rect 9890 24330 9920 24360
rect 10000 24330 10030 24360
rect 10230 24330 10260 24360
rect 10340 24330 10370 24360
rect 10620 24330 10650 24360
rect 10730 24330 10760 24360
rect 10880 24330 10910 24360
rect 10990 24330 11020 24360
rect 11220 24330 11250 24360
rect 11330 24330 11360 24360
rect 11620 24330 11650 24360
rect 11730 24330 11760 24360
rect 11880 24330 11910 24360
rect 11990 24330 12020 24360
rect 12220 24330 12250 24360
rect 12330 24330 12360 24360
rect 12600 24330 12630 24360
rect 12710 24330 12740 24360
rect 7430 23210 7460 23240
rect 7540 23210 7570 23240
rect 7690 23210 7720 23240
rect 7800 23210 7830 23240
rect 8030 23210 8060 23240
rect 8140 23210 8170 23240
rect 8550 23210 8580 23240
rect 8700 23210 8730 23240
rect 9290 23210 9320 23240
rect 9400 23210 9430 23240
rect 9630 23210 9660 23240
rect 9740 23210 9770 23240
rect 9890 23210 9920 23240
rect 10000 23210 10030 23240
rect 10230 23210 10260 23240
rect 10340 23210 10370 23240
rect 10620 23210 10650 23240
rect 10730 23210 10760 23240
rect 10880 23210 10910 23240
rect 10990 23210 11020 23240
rect 11220 23210 11250 23240
rect 11330 23210 11360 23240
rect 11620 23210 11650 23240
rect 11730 23210 11760 23240
rect 11880 23210 11910 23240
rect 11990 23210 12020 23240
rect 12220 23210 12250 23240
rect 12330 23210 12360 23240
rect 12600 23210 12630 23240
rect 12710 23210 12740 23240
rect 7430 22700 7460 22810
rect 7370 22680 7460 22700
rect 7370 22640 7380 22680
rect 7420 22640 7460 22680
rect 7370 22620 7460 22640
rect 7430 22570 7460 22620
rect 7540 22570 7570 22810
rect 7690 22790 7720 22810
rect 7630 22770 7720 22790
rect 7630 22730 7640 22770
rect 7680 22730 7720 22770
rect 7630 22710 7720 22730
rect 7430 22560 7570 22570
rect 7430 22520 7480 22560
rect 7520 22520 7570 22560
rect 7430 22510 7570 22520
rect 7690 22570 7720 22710
rect 7800 22570 7830 22810
rect 8030 22770 8060 23010
rect 8140 22770 8170 23010
rect 8930 22940 8960 22970
rect 8030 22740 8170 22770
rect 8030 22680 8060 22740
rect 7940 22670 8060 22680
rect 7940 22630 7960 22670
rect 8000 22630 8060 22670
rect 7940 22620 8060 22630
rect 7690 22560 7830 22570
rect 7690 22520 7740 22560
rect 7780 22520 7830 22560
rect 7690 22510 7830 22520
rect 7430 21700 7570 21710
rect 7430 21660 7480 21700
rect 7520 21660 7570 21700
rect 7430 21650 7570 21660
rect 7430 21580 7460 21650
rect 7540 21580 7570 21650
rect 7690 21680 7830 21690
rect 7690 21640 7740 21680
rect 7780 21640 7830 21680
rect 7690 21630 7830 21640
rect 7690 21580 7720 21630
rect 7800 21580 7830 21630
rect 8030 21580 8060 22620
rect 8140 21580 8170 22740
rect 8550 22690 8580 22810
rect 8700 22770 8730 22810
rect 8630 22750 8730 22770
rect 8630 22710 8650 22750
rect 8690 22710 8730 22750
rect 8630 22690 8730 22710
rect 8930 22690 8960 22740
rect 9290 22720 9320 23010
rect 8480 22670 8580 22690
rect 8480 22630 8500 22670
rect 8540 22630 8580 22670
rect 8480 22610 8580 22630
rect 8550 21570 8580 22610
rect 8700 21570 8730 22690
rect 8860 22670 8960 22690
rect 8860 22630 8880 22670
rect 8920 22630 8960 22670
rect 8860 22610 8960 22630
rect 9200 22700 9320 22720
rect 9200 22640 9220 22700
rect 9280 22640 9320 22700
rect 9200 22620 9320 22640
rect 8930 21570 8960 22610
rect 9290 21620 9320 22620
rect 9400 21620 9430 23010
rect 9630 22690 9660 22810
rect 9570 22670 9660 22690
rect 9570 22630 9580 22670
rect 9620 22630 9660 22670
rect 9570 22610 9660 22630
rect 9630 22560 9660 22610
rect 9740 22560 9770 22810
rect 9890 22790 9920 22810
rect 9830 22770 9920 22790
rect 9830 22730 9840 22770
rect 9880 22730 9920 22770
rect 9830 22710 9920 22730
rect 9630 22550 9770 22560
rect 9630 22510 9680 22550
rect 9720 22510 9770 22550
rect 9630 22500 9770 22510
rect 9890 22560 9920 22710
rect 10000 22560 10030 22810
rect 10230 22800 10260 23010
rect 10340 22800 10370 23010
rect 10230 22770 10370 22800
rect 10230 22670 10260 22770
rect 10140 22660 10260 22670
rect 10140 22620 10160 22660
rect 10200 22620 10260 22660
rect 10140 22610 10260 22620
rect 9890 22550 10030 22560
rect 9890 22510 9940 22550
rect 9980 22510 10030 22550
rect 9890 22500 10030 22510
rect 9290 21590 9430 21620
rect 9290 21570 9320 21590
rect 9400 21570 9430 21590
rect 9630 21670 9770 21680
rect 9630 21630 9680 21670
rect 9720 21630 9770 21670
rect 9630 21620 9770 21630
rect 9630 21570 9660 21620
rect 9740 21570 9770 21620
rect 9890 21670 10030 21680
rect 9890 21630 9940 21670
rect 9980 21630 10030 21670
rect 9890 21620 10030 21630
rect 9890 21570 9920 21620
rect 10000 21570 10030 21620
rect 10230 21570 10260 22610
rect 10340 21570 10370 22770
rect 10620 22690 10650 22810
rect 10560 22670 10650 22690
rect 10560 22630 10570 22670
rect 10610 22630 10650 22670
rect 10560 22610 10650 22630
rect 10620 22560 10650 22610
rect 10730 22560 10760 22810
rect 10880 22790 10910 22810
rect 10820 22770 10910 22790
rect 10820 22730 10830 22770
rect 10870 22730 10910 22770
rect 10820 22710 10910 22730
rect 10620 22550 10760 22560
rect 10620 22510 10670 22550
rect 10710 22510 10760 22550
rect 10620 22500 10760 22510
rect 10880 22560 10910 22710
rect 10990 22560 11020 22810
rect 11220 22770 11250 23010
rect 11330 22770 11360 23010
rect 12220 22810 12250 23010
rect 12330 22810 12360 23010
rect 11220 22740 11360 22770
rect 11220 22670 11250 22740
rect 11130 22660 11250 22670
rect 11130 22620 11150 22660
rect 11190 22620 11250 22660
rect 11130 22610 11250 22620
rect 10880 22550 11020 22560
rect 10880 22510 10930 22550
rect 10970 22510 11020 22550
rect 10880 22500 11020 22510
rect 10620 21670 10760 21680
rect 10620 21630 10670 21670
rect 10710 21630 10760 21670
rect 10620 21620 10760 21630
rect 10620 21570 10650 21620
rect 10730 21570 10760 21620
rect 10880 21670 11020 21680
rect 10880 21630 10930 21670
rect 10970 21630 11020 21670
rect 10880 21620 11020 21630
rect 10880 21570 10910 21620
rect 10990 21570 11020 21620
rect 11220 21570 11250 22610
rect 11330 21570 11360 22740
rect 11620 22690 11650 22810
rect 11560 22670 11650 22690
rect 11560 22630 11570 22670
rect 11610 22630 11650 22670
rect 11560 22610 11650 22630
rect 11620 22560 11650 22610
rect 11730 22560 11760 22810
rect 11880 22790 11910 22810
rect 11820 22770 11910 22790
rect 11820 22730 11830 22770
rect 11870 22730 11910 22770
rect 11820 22710 11910 22730
rect 11620 22550 11760 22560
rect 11620 22510 11670 22550
rect 11710 22510 11760 22550
rect 11620 22500 11760 22510
rect 11880 22560 11910 22710
rect 11990 22560 12020 22810
rect 12220 22780 12360 22810
rect 12220 22670 12250 22780
rect 12130 22660 12250 22670
rect 12130 22620 12150 22660
rect 12190 22620 12250 22660
rect 12130 22610 12250 22620
rect 11880 22550 12020 22560
rect 11880 22510 11930 22550
rect 11970 22510 12020 22550
rect 11880 22500 12020 22510
rect 11620 21670 11760 21680
rect 11620 21630 11670 21670
rect 11710 21630 11760 21670
rect 11620 21620 11760 21630
rect 11620 21570 11650 21620
rect 11730 21570 11760 21620
rect 11880 21670 12020 21680
rect 11880 21630 11930 21670
rect 11970 21630 12020 21670
rect 11880 21620 12020 21630
rect 11880 21570 11910 21620
rect 11990 21570 12020 21620
rect 12220 21570 12250 22610
rect 12330 21570 12360 22780
rect 12600 22820 12630 23010
rect 12710 22820 12740 23010
rect 12950 22930 12980 22960
rect 13180 22930 13210 22960
rect 13290 22930 13320 22960
rect 13520 22930 13550 22960
rect 13630 22930 13660 22960
rect 13740 22930 13770 22960
rect 13850 22930 13880 22960
rect 14080 22930 14110 22960
rect 14190 22930 14220 22960
rect 14300 22930 14330 22960
rect 14410 22930 14440 22960
rect 14520 22930 14550 22960
rect 14630 22930 14660 22960
rect 14740 22930 14770 22960
rect 14850 22930 14880 22960
rect 15140 22930 15170 22960
rect 15250 22930 15280 22960
rect 15360 22930 15390 22960
rect 15470 22930 15500 22960
rect 15580 22930 15610 22960
rect 15690 22930 15720 22960
rect 15800 22930 15830 22960
rect 15910 22930 15940 22960
rect 16020 22930 16050 22960
rect 16130 22930 16160 22960
rect 16240 22930 16270 22960
rect 16350 22930 16380 22960
rect 16460 22930 16490 22960
rect 16570 22930 16600 22960
rect 16680 22930 16710 22960
rect 16790 22930 16820 22960
rect 17090 22930 17120 22960
rect 17200 22930 17230 22960
rect 17310 22930 17340 22960
rect 17420 22930 17450 22960
rect 17530 22930 17560 22960
rect 17640 22930 17670 22960
rect 17750 22930 17780 22960
rect 17860 22930 17890 22960
rect 17970 22930 18000 22960
rect 18080 22930 18110 22960
rect 18190 22930 18220 22960
rect 18300 22930 18330 22960
rect 18410 22930 18440 22960
rect 18520 22930 18550 22960
rect 18630 22930 18660 22960
rect 18740 22930 18770 22960
rect 18850 22930 18880 22960
rect 18960 22930 18990 22960
rect 19070 22930 19100 22960
rect 19180 22930 19210 22960
rect 19290 22930 19320 22960
rect 19400 22930 19430 22960
rect 19510 22930 19540 22960
rect 19620 22930 19650 22960
rect 19730 22930 19760 22960
rect 19840 22930 19870 22960
rect 19950 22930 19980 22960
rect 20060 22930 20090 22960
rect 20170 22930 20200 22960
rect 20280 22930 20310 22960
rect 20390 22930 20420 22960
rect 20500 22930 20530 22960
rect 12600 22790 12740 22820
rect 12600 22670 12630 22790
rect 12510 22660 12630 22670
rect 12510 22620 12530 22660
rect 12570 22620 12630 22660
rect 12510 22610 12630 22620
rect 12600 21570 12630 22610
rect 12710 21570 12740 22790
rect 12950 22690 12980 22730
rect 13180 22690 13210 22730
rect 13290 22690 13320 22730
rect 13520 22690 13550 22730
rect 13630 22690 13660 22730
rect 13740 22690 13770 22730
rect 13850 22690 13880 22730
rect 14080 22690 14110 22730
rect 14190 22690 14220 22730
rect 14300 22690 14330 22730
rect 14410 22690 14440 22730
rect 14520 22690 14550 22730
rect 14630 22690 14660 22730
rect 14740 22690 14770 22730
rect 14850 22690 14880 22730
rect 15140 22690 15170 22730
rect 15250 22690 15280 22730
rect 15360 22690 15390 22730
rect 15470 22690 15500 22730
rect 15580 22690 15610 22730
rect 15690 22690 15720 22730
rect 15800 22690 15830 22730
rect 15910 22690 15940 22730
rect 16020 22690 16050 22730
rect 16130 22690 16160 22730
rect 16240 22690 16270 22730
rect 16350 22690 16380 22730
rect 16460 22690 16490 22730
rect 16570 22690 16600 22730
rect 16680 22690 16710 22730
rect 16790 22690 16820 22730
rect 17090 22690 17120 22730
rect 17200 22690 17230 22730
rect 17310 22690 17340 22730
rect 17420 22690 17450 22730
rect 17530 22690 17560 22730
rect 17640 22690 17670 22730
rect 17750 22690 17780 22730
rect 17860 22690 17890 22730
rect 17970 22690 18000 22730
rect 18080 22690 18110 22730
rect 18190 22690 18220 22730
rect 18300 22690 18330 22730
rect 18410 22690 18440 22730
rect 18520 22690 18550 22730
rect 18630 22690 18660 22730
rect 18740 22690 18770 22730
rect 18850 22690 18880 22730
rect 18960 22690 18990 22730
rect 19070 22690 19100 22730
rect 19180 22690 19210 22730
rect 19290 22690 19320 22730
rect 19400 22690 19430 22730
rect 19510 22690 19540 22730
rect 19620 22690 19650 22730
rect 19730 22690 19760 22730
rect 19840 22690 19870 22730
rect 19950 22690 19980 22730
rect 20060 22690 20090 22730
rect 20170 22690 20200 22730
rect 20280 22690 20310 22730
rect 20390 22690 20420 22730
rect 20500 22690 20530 22730
rect 12890 22670 12980 22690
rect 12890 22630 12900 22670
rect 12940 22630 12980 22670
rect 12890 22610 12980 22630
rect 13120 22670 13320 22690
rect 13120 22630 13130 22670
rect 13170 22650 13320 22670
rect 13170 22630 13210 22650
rect 13120 22610 13210 22630
rect 12950 21570 12980 22610
rect 13180 22580 13210 22610
rect 13290 22580 13320 22650
rect 13460 22670 13880 22690
rect 13460 22630 13470 22670
rect 13510 22650 13880 22670
rect 13510 22630 13550 22650
rect 13460 22610 13550 22630
rect 13180 22570 13320 22580
rect 13180 22530 13230 22570
rect 13270 22530 13320 22570
rect 13180 22520 13320 22530
rect 13520 22580 13550 22610
rect 13630 22580 13660 22650
rect 13520 22570 13660 22580
rect 13520 22530 13570 22570
rect 13610 22530 13660 22570
rect 13520 22520 13660 22530
rect 13740 22580 13770 22650
rect 13850 22580 13880 22650
rect 14020 22670 14880 22690
rect 14020 22630 14030 22670
rect 14070 22650 14880 22670
rect 14070 22630 14110 22650
rect 14020 22610 14110 22630
rect 13740 22570 13880 22580
rect 13740 22530 13790 22570
rect 13830 22530 13880 22570
rect 13740 22520 13880 22530
rect 14080 22560 14110 22610
rect 14190 22560 14220 22650
rect 14080 22550 14220 22560
rect 14080 22510 14130 22550
rect 14170 22510 14220 22550
rect 14080 22500 14220 22510
rect 14300 22560 14330 22650
rect 14410 22560 14440 22650
rect 14300 22550 14440 22560
rect 14300 22510 14350 22550
rect 14390 22510 14440 22550
rect 14300 22500 14440 22510
rect 14520 22560 14550 22650
rect 14630 22560 14660 22650
rect 14520 22550 14660 22560
rect 14520 22510 14570 22550
rect 14610 22510 14660 22550
rect 14520 22500 14660 22510
rect 14740 22560 14770 22650
rect 14850 22560 14880 22650
rect 15080 22670 16820 22690
rect 15080 22630 15090 22670
rect 15130 22650 16820 22670
rect 15130 22630 15170 22650
rect 15080 22610 15170 22630
rect 14740 22550 14880 22560
rect 14740 22510 14790 22550
rect 14830 22510 14880 22550
rect 14740 22500 14880 22510
rect 15140 22560 15170 22610
rect 15250 22560 15280 22650
rect 15140 22550 15280 22560
rect 15140 22510 15190 22550
rect 15230 22510 15280 22550
rect 15140 22500 15280 22510
rect 15360 22560 15390 22650
rect 15470 22560 15500 22650
rect 15360 22550 15500 22560
rect 15360 22510 15410 22550
rect 15450 22510 15500 22550
rect 15360 22500 15500 22510
rect 15580 22560 15610 22650
rect 15690 22560 15720 22650
rect 15580 22550 15720 22560
rect 15580 22510 15630 22550
rect 15670 22510 15720 22550
rect 15580 22500 15720 22510
rect 15800 22560 15830 22650
rect 15910 22560 15940 22650
rect 15800 22550 15940 22560
rect 15800 22510 15850 22550
rect 15890 22510 15940 22550
rect 15800 22500 15940 22510
rect 16020 22560 16050 22650
rect 16130 22560 16160 22650
rect 16020 22550 16160 22560
rect 16020 22510 16070 22550
rect 16110 22510 16160 22550
rect 16020 22500 16160 22510
rect 16240 22560 16270 22650
rect 16350 22560 16380 22650
rect 16240 22550 16380 22560
rect 16240 22510 16290 22550
rect 16330 22510 16380 22550
rect 16240 22500 16380 22510
rect 16460 22560 16490 22650
rect 16570 22560 16600 22650
rect 16460 22550 16600 22560
rect 16460 22510 16510 22550
rect 16550 22510 16600 22550
rect 16460 22500 16600 22510
rect 16680 22560 16710 22650
rect 16790 22560 16820 22650
rect 17020 22670 20530 22690
rect 17020 22630 17040 22670
rect 17080 22650 20530 22670
rect 17080 22630 17120 22650
rect 17020 22610 17120 22630
rect 16680 22550 16820 22560
rect 16680 22510 16730 22550
rect 16770 22510 16820 22550
rect 16680 22500 16820 22510
rect 17090 22560 17120 22610
rect 17200 22560 17230 22650
rect 17090 22550 17230 22560
rect 17090 22510 17140 22550
rect 17180 22510 17230 22550
rect 17090 22500 17230 22510
rect 17310 22560 17340 22650
rect 17420 22560 17450 22650
rect 17310 22550 17450 22560
rect 17310 22510 17360 22550
rect 17400 22510 17450 22550
rect 17310 22500 17450 22510
rect 17530 22560 17560 22650
rect 17640 22560 17670 22650
rect 17530 22550 17670 22560
rect 17530 22510 17580 22550
rect 17620 22510 17670 22550
rect 17530 22500 17670 22510
rect 17750 22560 17780 22650
rect 17860 22560 17890 22650
rect 17750 22550 17890 22560
rect 17750 22510 17800 22550
rect 17840 22510 17890 22550
rect 17750 22500 17890 22510
rect 17970 22560 18000 22650
rect 18080 22560 18110 22650
rect 17970 22550 18110 22560
rect 17970 22510 18020 22550
rect 18060 22510 18110 22550
rect 17970 22500 18110 22510
rect 18190 22560 18220 22650
rect 18300 22560 18330 22650
rect 18190 22550 18330 22560
rect 18190 22510 18240 22550
rect 18280 22510 18330 22550
rect 18190 22500 18330 22510
rect 18410 22560 18440 22650
rect 18520 22560 18550 22650
rect 18410 22550 18550 22560
rect 18410 22510 18460 22550
rect 18500 22510 18550 22550
rect 18410 22500 18550 22510
rect 18630 22560 18660 22650
rect 18740 22560 18770 22650
rect 18630 22550 18770 22560
rect 18630 22510 18680 22550
rect 18720 22510 18770 22550
rect 18630 22500 18770 22510
rect 18850 22560 18880 22650
rect 18960 22560 18990 22650
rect 18850 22550 18990 22560
rect 18850 22510 18900 22550
rect 18940 22510 18990 22550
rect 18850 22500 18990 22510
rect 19070 22560 19100 22650
rect 19180 22560 19210 22650
rect 19070 22550 19210 22560
rect 19070 22510 19120 22550
rect 19160 22510 19210 22550
rect 19070 22500 19210 22510
rect 19290 22560 19320 22650
rect 19400 22560 19430 22650
rect 19290 22550 19430 22560
rect 19290 22510 19340 22550
rect 19380 22510 19430 22550
rect 19290 22500 19430 22510
rect 19510 22560 19540 22650
rect 19620 22560 19650 22650
rect 19510 22550 19650 22560
rect 19510 22510 19560 22550
rect 19600 22510 19650 22550
rect 19510 22500 19650 22510
rect 19730 22560 19760 22650
rect 19840 22560 19870 22650
rect 19730 22550 19870 22560
rect 19730 22510 19780 22550
rect 19820 22510 19870 22550
rect 19730 22500 19870 22510
rect 19950 22560 19980 22650
rect 20060 22560 20090 22650
rect 19950 22550 20090 22560
rect 19950 22510 20000 22550
rect 20040 22510 20090 22550
rect 19950 22500 20090 22510
rect 20170 22560 20200 22650
rect 20280 22560 20310 22650
rect 20170 22550 20310 22560
rect 20170 22510 20220 22550
rect 20260 22510 20310 22550
rect 20170 22500 20310 22510
rect 20390 22560 20420 22650
rect 20500 22560 20530 22650
rect 20390 22550 20530 22560
rect 20390 22510 20440 22550
rect 20480 22510 20530 22550
rect 20390 22500 20530 22510
rect 13180 21680 13320 21690
rect 13180 21640 13230 21680
rect 13270 21640 13320 21680
rect 13180 21630 13320 21640
rect 13180 21570 13210 21630
rect 13290 21570 13320 21630
rect 13520 21680 13660 21690
rect 13520 21640 13570 21680
rect 13610 21640 13660 21680
rect 13520 21630 13660 21640
rect 13520 21570 13550 21630
rect 13630 21570 13660 21630
rect 13740 21680 13880 21690
rect 13740 21640 13790 21680
rect 13830 21640 13880 21680
rect 13740 21630 13880 21640
rect 13740 21570 13770 21630
rect 13850 21570 13880 21630
rect 14080 21660 14220 21670
rect 14080 21620 14130 21660
rect 14170 21620 14220 21660
rect 14080 21610 14220 21620
rect 14080 21570 14110 21610
rect 14190 21570 14220 21610
rect 14300 21660 14440 21670
rect 14300 21620 14350 21660
rect 14390 21620 14440 21660
rect 14300 21610 14440 21620
rect 14300 21570 14330 21610
rect 14410 21570 14440 21610
rect 14520 21660 14660 21670
rect 14520 21620 14570 21660
rect 14610 21620 14660 21660
rect 14520 21610 14660 21620
rect 14520 21570 14550 21610
rect 14630 21570 14660 21610
rect 14740 21660 14880 21670
rect 14740 21620 14790 21660
rect 14830 21620 14880 21660
rect 14740 21610 14880 21620
rect 14740 21570 14770 21610
rect 14850 21570 14880 21610
rect 15140 21660 15280 21670
rect 15140 21620 15190 21660
rect 15230 21620 15280 21660
rect 15140 21610 15280 21620
rect 15140 21570 15170 21610
rect 15250 21570 15280 21610
rect 15360 21660 15500 21670
rect 15360 21620 15410 21660
rect 15450 21620 15500 21660
rect 15360 21610 15500 21620
rect 15360 21570 15390 21610
rect 15470 21570 15500 21610
rect 15580 21660 15720 21670
rect 15580 21620 15630 21660
rect 15670 21620 15720 21660
rect 15580 21610 15720 21620
rect 15580 21570 15610 21610
rect 15690 21570 15720 21610
rect 15800 21660 15940 21670
rect 15800 21620 15850 21660
rect 15890 21620 15940 21660
rect 15800 21610 15940 21620
rect 15800 21570 15830 21610
rect 15910 21570 15940 21610
rect 16020 21660 16160 21670
rect 16020 21620 16070 21660
rect 16110 21620 16160 21660
rect 16020 21610 16160 21620
rect 16020 21570 16050 21610
rect 16130 21570 16160 21610
rect 16240 21660 16380 21670
rect 16240 21620 16290 21660
rect 16330 21620 16380 21660
rect 16240 21610 16380 21620
rect 16240 21570 16270 21610
rect 16350 21570 16380 21610
rect 16460 21660 16600 21670
rect 16460 21620 16510 21660
rect 16550 21620 16600 21660
rect 16460 21610 16600 21620
rect 16460 21570 16490 21610
rect 16570 21570 16600 21610
rect 16680 21660 16820 21670
rect 16680 21620 16730 21660
rect 16770 21620 16820 21660
rect 16680 21610 16820 21620
rect 16680 21570 16710 21610
rect 16790 21570 16820 21610
rect 17090 21660 17230 21670
rect 17090 21620 17140 21660
rect 17180 21620 17230 21660
rect 17090 21610 17230 21620
rect 17090 21570 17120 21610
rect 17200 21570 17230 21610
rect 17310 21660 17450 21670
rect 17310 21620 17360 21660
rect 17400 21620 17450 21660
rect 17310 21610 17450 21620
rect 17310 21570 17340 21610
rect 17420 21570 17450 21610
rect 17530 21660 17670 21670
rect 17530 21620 17580 21660
rect 17620 21620 17670 21660
rect 17530 21610 17670 21620
rect 17530 21570 17560 21610
rect 17640 21570 17670 21610
rect 17750 21660 17890 21670
rect 17750 21620 17800 21660
rect 17840 21620 17890 21660
rect 17750 21610 17890 21620
rect 17750 21570 17780 21610
rect 17860 21570 17890 21610
rect 17970 21660 18110 21670
rect 17970 21620 18020 21660
rect 18060 21620 18110 21660
rect 17970 21610 18110 21620
rect 17970 21570 18000 21610
rect 18080 21570 18110 21610
rect 18190 21660 18330 21670
rect 18190 21620 18240 21660
rect 18280 21620 18330 21660
rect 18190 21610 18330 21620
rect 18190 21570 18220 21610
rect 18300 21570 18330 21610
rect 18410 21660 18550 21670
rect 18410 21620 18460 21660
rect 18500 21620 18550 21660
rect 18410 21610 18550 21620
rect 18410 21570 18440 21610
rect 18520 21570 18550 21610
rect 18630 21660 18770 21670
rect 18630 21620 18680 21660
rect 18720 21620 18770 21660
rect 18630 21610 18770 21620
rect 18630 21570 18660 21610
rect 18740 21570 18770 21610
rect 18850 21660 18990 21670
rect 18850 21620 18900 21660
rect 18940 21620 18990 21660
rect 18850 21610 18990 21620
rect 18850 21570 18880 21610
rect 18960 21570 18990 21610
rect 19070 21660 19210 21670
rect 19070 21620 19120 21660
rect 19160 21620 19210 21660
rect 19070 21610 19210 21620
rect 19070 21570 19100 21610
rect 19180 21570 19210 21610
rect 19290 21660 19430 21670
rect 19290 21620 19340 21660
rect 19380 21620 19430 21660
rect 19290 21610 19430 21620
rect 19290 21570 19320 21610
rect 19400 21570 19430 21610
rect 19510 21660 19650 21670
rect 19510 21620 19560 21660
rect 19600 21620 19650 21660
rect 19510 21610 19650 21620
rect 19510 21570 19540 21610
rect 19620 21570 19650 21610
rect 19730 21660 19870 21670
rect 19730 21620 19780 21660
rect 19820 21620 19870 21660
rect 19730 21610 19870 21620
rect 19730 21570 19760 21610
rect 19840 21570 19870 21610
rect 19950 21660 20090 21670
rect 19950 21620 20000 21660
rect 20040 21620 20090 21660
rect 19950 21610 20090 21620
rect 19950 21570 19980 21610
rect 20060 21570 20090 21610
rect 20170 21660 20310 21670
rect 20170 21620 20220 21660
rect 20260 21620 20310 21660
rect 20170 21610 20310 21620
rect 20170 21570 20200 21610
rect 20280 21570 20310 21610
rect 20390 21660 20530 21670
rect 20390 21620 20440 21660
rect 20480 21620 20530 21660
rect 20390 21610 20530 21620
rect 20390 21570 20420 21610
rect 20500 21570 20530 21610
rect 7430 21050 7460 21080
rect 7540 21050 7570 21080
rect 7690 21050 7720 21080
rect 7800 21050 7830 21080
rect 8030 21050 8060 21080
rect 8140 21050 8170 21080
rect 8550 21040 8580 21070
rect 8700 21040 8730 21070
rect 8930 21040 8960 21070
rect 9290 21040 9320 21070
rect 9400 21040 9430 21070
rect 9630 21040 9660 21070
rect 9740 21040 9770 21070
rect 9890 21040 9920 21070
rect 10000 21040 10030 21070
rect 10230 21040 10260 21070
rect 10340 21040 10370 21070
rect 10620 21040 10650 21070
rect 10730 21040 10760 21070
rect 10880 21040 10910 21070
rect 10990 21040 11020 21070
rect 11220 21040 11250 21070
rect 11330 21040 11360 21070
rect 11620 21040 11650 21070
rect 11730 21040 11760 21070
rect 11880 21040 11910 21070
rect 11990 21040 12020 21070
rect 12220 21040 12250 21070
rect 12330 21040 12360 21070
rect 12600 21040 12630 21070
rect 12710 21040 12740 21070
rect 12950 21040 12980 21070
rect 13180 21040 13210 21070
rect 13290 21040 13320 21070
rect 13520 21040 13550 21070
rect 13630 21040 13660 21070
rect 13740 21040 13770 21070
rect 13850 21040 13880 21070
rect 14080 21040 14110 21070
rect 14190 21040 14220 21070
rect 14300 21040 14330 21070
rect 14410 21040 14440 21070
rect 14520 21040 14550 21070
rect 14630 21040 14660 21070
rect 14740 21040 14770 21070
rect 14850 21040 14880 21070
rect 15140 21040 15170 21070
rect 15250 21040 15280 21070
rect 15360 21040 15390 21070
rect 15470 21040 15500 21070
rect 15580 21040 15610 21070
rect 15690 21040 15720 21070
rect 15800 21040 15830 21070
rect 15910 21040 15940 21070
rect 16020 21040 16050 21070
rect 16130 21040 16160 21070
rect 16240 21040 16270 21070
rect 16350 21040 16380 21070
rect 16460 21040 16490 21070
rect 16570 21040 16600 21070
rect 16680 21040 16710 21070
rect 16790 21040 16820 21070
rect 17090 21040 17120 21070
rect 17200 21040 17230 21070
rect 17310 21040 17340 21070
rect 17420 21040 17450 21070
rect 17530 21040 17560 21070
rect 17640 21040 17670 21070
rect 17750 21040 17780 21070
rect 17860 21040 17890 21070
rect 17970 21040 18000 21070
rect 18080 21040 18110 21070
rect 18190 21040 18220 21070
rect 18300 21040 18330 21070
rect 18410 21040 18440 21070
rect 18520 21040 18550 21070
rect 18630 21040 18660 21070
rect 18740 21040 18770 21070
rect 18850 21040 18880 21070
rect 18960 21040 18990 21070
rect 19070 21040 19100 21070
rect 19180 21040 19210 21070
rect 19290 21040 19320 21070
rect 19400 21040 19430 21070
rect 19510 21040 19540 21070
rect 19620 21040 19650 21070
rect 19730 21040 19760 21070
rect 19840 21040 19870 21070
rect 19950 21040 19980 21070
rect 20060 21040 20090 21070
rect 20170 21040 20200 21070
rect 20280 21040 20310 21070
rect 20390 21040 20420 21070
rect 20500 21040 20530 21070
rect 7350 20360 7380 20390
rect 7460 20360 7490 20390
rect 7610 20360 7640 20390
rect 7720 20360 7750 20390
rect 8020 20360 8050 20390
rect 8130 20360 8160 20390
rect 8550 19910 8580 19940
rect 8700 19910 8730 19940
rect 8930 19910 8960 19940
rect 9290 19910 9320 19940
rect 9400 19910 9430 19940
rect 9630 19910 9660 19940
rect 9740 19910 9770 19940
rect 9890 19910 9920 19940
rect 10000 19910 10030 19940
rect 10230 19910 10260 19940
rect 10340 19910 10370 19940
rect 10620 19910 10650 19940
rect 10730 19910 10760 19940
rect 10880 19910 10910 19940
rect 10990 19910 11020 19940
rect 11220 19910 11250 19940
rect 11330 19910 11360 19940
rect 11620 19910 11650 19940
rect 11730 19910 11760 19940
rect 11880 19910 11910 19940
rect 11990 19910 12020 19940
rect 12220 19910 12250 19940
rect 12330 19910 12360 19940
rect 12600 19910 12630 19940
rect 12710 19910 12740 19940
rect 12950 19910 12980 19940
rect 13180 19910 13210 19940
rect 13290 19910 13320 19940
rect 13520 19910 13550 19940
rect 13630 19910 13660 19940
rect 13740 19910 13770 19940
rect 13850 19910 13880 19940
rect 14080 19910 14110 19940
rect 14190 19910 14220 19940
rect 14300 19910 14330 19940
rect 14410 19910 14440 19940
rect 14520 19910 14550 19940
rect 14630 19910 14660 19940
rect 14740 19910 14770 19940
rect 14850 19910 14880 19940
rect 15140 19910 15170 19940
rect 15250 19910 15280 19940
rect 15360 19910 15390 19940
rect 15470 19910 15500 19940
rect 15580 19910 15610 19940
rect 15690 19910 15720 19940
rect 15800 19910 15830 19940
rect 15910 19910 15940 19940
rect 16020 19910 16050 19940
rect 16130 19910 16160 19940
rect 16240 19910 16270 19940
rect 16350 19910 16380 19940
rect 16460 19910 16490 19940
rect 16570 19910 16600 19940
rect 16680 19910 16710 19940
rect 16790 19910 16820 19940
rect 17090 19910 17120 19940
rect 17200 19910 17230 19940
rect 17310 19910 17340 19940
rect 17420 19910 17450 19940
rect 17530 19910 17560 19940
rect 17640 19910 17670 19940
rect 17750 19910 17780 19940
rect 17860 19910 17890 19940
rect 17970 19910 18000 19940
rect 18080 19910 18110 19940
rect 18190 19910 18220 19940
rect 18300 19910 18330 19940
rect 18410 19910 18440 19940
rect 18520 19910 18550 19940
rect 18630 19910 18660 19940
rect 18740 19910 18770 19940
rect 18850 19910 18880 19940
rect 18960 19910 18990 19940
rect 19070 19910 19100 19940
rect 19180 19910 19210 19940
rect 19290 19910 19320 19940
rect 19400 19910 19430 19940
rect 19510 19910 19540 19940
rect 19620 19910 19650 19940
rect 19730 19910 19760 19940
rect 19840 19910 19870 19940
rect 19950 19910 19980 19940
rect 20060 19910 20090 19940
rect 20170 19910 20200 19940
rect 20280 19910 20310 19940
rect 20390 19910 20420 19940
rect 20500 19910 20530 19940
rect 7350 19320 7380 19360
rect 7460 19320 7490 19360
rect 7350 19310 7490 19320
rect 7350 19270 7400 19310
rect 7440 19270 7490 19310
rect 7350 19260 7490 19270
rect 7350 18430 7490 18440
rect 7350 18390 7400 18430
rect 7440 18390 7490 18430
rect 7350 18380 7490 18390
rect 7350 18190 7380 18380
rect 7290 18170 7380 18190
rect 7290 18130 7300 18170
rect 7340 18130 7380 18170
rect 7290 18110 7380 18130
rect 7350 17980 7380 18110
rect 7460 17980 7490 18380
rect 7610 18300 7640 19360
rect 7550 18280 7640 18300
rect 7720 18280 7750 19360
rect 8020 18300 8050 19860
rect 7550 18240 7560 18280
rect 7600 18250 7750 18280
rect 7600 18240 7640 18250
rect 7550 18220 7640 18240
rect 7610 17980 7640 18220
rect 7720 17980 7750 18250
rect 7960 18280 8050 18300
rect 7960 18240 7970 18280
rect 8010 18270 8050 18280
rect 8130 18270 8160 19860
rect 8550 18370 8580 19410
rect 8480 18350 8580 18370
rect 8480 18310 8500 18350
rect 8540 18310 8580 18350
rect 8480 18290 8580 18310
rect 8700 18290 8730 19410
rect 8930 18370 8960 19410
rect 8860 18350 8960 18370
rect 9290 18350 9320 19410
rect 8860 18310 8880 18350
rect 8920 18310 8960 18350
rect 8860 18290 8960 18310
rect 8010 18240 8160 18270
rect 7960 18220 8050 18240
rect 8020 17980 8050 18220
rect 8130 17980 8160 18240
rect 8550 18170 8580 18290
rect 8630 18270 8730 18290
rect 8630 18230 8650 18270
rect 8690 18230 8730 18270
rect 8930 18240 8960 18290
rect 9200 18330 9320 18350
rect 9200 18270 9220 18330
rect 9280 18320 9320 18330
rect 9400 18320 9430 19410
rect 9630 19370 9660 19410
rect 9740 19370 9770 19410
rect 9630 19360 9770 19370
rect 9630 19320 9680 19360
rect 9720 19320 9770 19360
rect 9630 19310 9770 19320
rect 9890 19370 9920 19410
rect 10000 19370 10030 19410
rect 9890 19360 10030 19370
rect 9890 19320 9940 19360
rect 9980 19320 10030 19360
rect 9890 19310 10030 19320
rect 9630 18470 9770 18480
rect 9630 18430 9680 18470
rect 9720 18430 9770 18470
rect 9630 18420 9770 18430
rect 9630 18370 9660 18420
rect 9280 18280 9430 18320
rect 9570 18350 9660 18370
rect 9570 18310 9580 18350
rect 9620 18310 9660 18350
rect 9570 18290 9660 18310
rect 9280 18270 9320 18280
rect 9200 18250 9320 18270
rect 8630 18210 8730 18230
rect 8700 18170 8730 18210
rect 7350 17740 7380 17780
rect 7460 17740 7490 17780
rect 7610 17740 7640 17780
rect 7720 17740 7750 17780
rect 8020 17740 8050 17780
rect 8130 17740 8160 17780
rect 8930 18010 8960 18040
rect 9290 17970 9320 18250
rect 9400 17970 9430 18280
rect 9630 18170 9660 18290
rect 9740 18170 9770 18420
rect 9890 18470 10030 18480
rect 9890 18430 9940 18470
rect 9980 18430 10030 18470
rect 9890 18420 10030 18430
rect 9890 18270 9920 18420
rect 9830 18250 9920 18270
rect 9830 18210 9840 18250
rect 9880 18210 9920 18250
rect 9830 18190 9920 18210
rect 9890 18170 9920 18190
rect 10000 18170 10030 18420
rect 10230 18370 10260 19410
rect 10140 18360 10260 18370
rect 10140 18320 10160 18360
rect 10200 18320 10260 18360
rect 10140 18310 10260 18320
rect 10230 18290 10260 18310
rect 10340 18290 10370 19410
rect 10620 19370 10650 19410
rect 10730 19370 10760 19410
rect 10620 19360 10760 19370
rect 10620 19320 10670 19360
rect 10710 19320 10760 19360
rect 10620 19310 10760 19320
rect 10880 19370 10910 19410
rect 10990 19370 11020 19410
rect 10880 19360 11020 19370
rect 10880 19320 10930 19360
rect 10970 19320 11020 19360
rect 10880 19310 11020 19320
rect 10620 18470 10760 18480
rect 10620 18430 10670 18470
rect 10710 18430 10760 18470
rect 10620 18420 10760 18430
rect 10620 18370 10650 18420
rect 10560 18350 10650 18370
rect 10560 18310 10570 18350
rect 10610 18310 10650 18350
rect 10560 18290 10650 18310
rect 10230 18260 10370 18290
rect 10230 17970 10260 18260
rect 10340 17970 10370 18260
rect 10620 18170 10650 18290
rect 10730 18170 10760 18420
rect 10880 18470 11020 18480
rect 10880 18430 10930 18470
rect 10970 18430 11020 18470
rect 10880 18420 11020 18430
rect 10880 18270 10910 18420
rect 10820 18250 10910 18270
rect 10820 18210 10830 18250
rect 10870 18210 10910 18250
rect 10820 18190 10910 18210
rect 10880 18170 10910 18190
rect 10990 18170 11020 18420
rect 11220 18370 11250 19410
rect 11130 18360 11250 18370
rect 11130 18320 11150 18360
rect 11190 18320 11250 18360
rect 11130 18310 11250 18320
rect 11220 18290 11250 18310
rect 11330 18290 11360 19410
rect 11620 19360 11650 19410
rect 11730 19360 11760 19410
rect 11620 19350 11760 19360
rect 11620 19310 11670 19350
rect 11710 19310 11760 19350
rect 11620 19300 11760 19310
rect 11880 19360 11910 19410
rect 11990 19360 12020 19410
rect 11880 19350 12020 19360
rect 11880 19310 11930 19350
rect 11970 19310 12020 19350
rect 11880 19300 12020 19310
rect 11620 18460 11760 18470
rect 11620 18420 11670 18460
rect 11710 18420 11760 18460
rect 11620 18410 11760 18420
rect 11620 18370 11650 18410
rect 11560 18350 11650 18370
rect 11560 18310 11570 18350
rect 11610 18310 11650 18350
rect 11560 18290 11650 18310
rect 11220 18260 11360 18290
rect 11220 17970 11250 18260
rect 11330 17970 11360 18260
rect 11620 18170 11650 18290
rect 11730 18170 11760 18410
rect 11880 18460 12020 18470
rect 11880 18420 11930 18460
rect 11970 18420 12020 18460
rect 11880 18410 12020 18420
rect 11880 18270 11910 18410
rect 11820 18250 11910 18270
rect 11820 18210 11830 18250
rect 11870 18210 11910 18250
rect 11820 18190 11910 18210
rect 11880 18170 11910 18190
rect 11990 18170 12020 18410
rect 12220 18370 12250 19410
rect 12130 18360 12250 18370
rect 12130 18320 12150 18360
rect 12190 18320 12250 18360
rect 12130 18310 12250 18320
rect 12220 18300 12250 18310
rect 12330 18300 12360 19410
rect 12600 18370 12630 19410
rect 12510 18360 12630 18370
rect 12510 18320 12530 18360
rect 12570 18320 12630 18360
rect 12510 18310 12630 18320
rect 12220 18270 12360 18300
rect 12220 17970 12250 18270
rect 12330 17970 12360 18270
rect 12600 18250 12630 18310
rect 12710 18250 12740 19410
rect 12950 18370 12980 19410
rect 13180 19350 13210 19410
rect 13290 19350 13320 19410
rect 13180 19340 13320 19350
rect 13180 19300 13230 19340
rect 13270 19300 13320 19340
rect 13180 19290 13320 19300
rect 13520 19350 13550 19410
rect 13630 19350 13660 19410
rect 13520 19340 13660 19350
rect 13520 19300 13570 19340
rect 13610 19300 13660 19340
rect 13520 19290 13660 19300
rect 13740 19350 13770 19410
rect 13850 19350 13880 19410
rect 13740 19340 13880 19350
rect 13740 19300 13790 19340
rect 13830 19300 13880 19340
rect 14080 19370 14110 19410
rect 14190 19370 14220 19410
rect 14080 19360 14220 19370
rect 14080 19320 14130 19360
rect 14170 19320 14220 19360
rect 14080 19310 14220 19320
rect 14300 19370 14330 19410
rect 14410 19370 14440 19410
rect 14300 19360 14440 19370
rect 14300 19320 14350 19360
rect 14390 19320 14440 19360
rect 14300 19310 14440 19320
rect 14520 19370 14550 19410
rect 14630 19370 14660 19410
rect 14520 19360 14660 19370
rect 14520 19320 14570 19360
rect 14610 19320 14660 19360
rect 14520 19310 14660 19320
rect 14740 19370 14770 19410
rect 14850 19370 14880 19410
rect 14740 19360 14880 19370
rect 14740 19320 14790 19360
rect 14830 19320 14880 19360
rect 14740 19310 14880 19320
rect 15140 19370 15170 19410
rect 15250 19370 15280 19410
rect 15140 19360 15280 19370
rect 15140 19320 15190 19360
rect 15230 19320 15280 19360
rect 15140 19310 15280 19320
rect 15360 19370 15390 19410
rect 15470 19370 15500 19410
rect 15360 19360 15500 19370
rect 15360 19320 15410 19360
rect 15450 19320 15500 19360
rect 15360 19310 15500 19320
rect 15580 19370 15610 19410
rect 15690 19370 15720 19410
rect 15580 19360 15720 19370
rect 15580 19320 15630 19360
rect 15670 19320 15720 19360
rect 15580 19310 15720 19320
rect 15800 19370 15830 19410
rect 15910 19370 15940 19410
rect 15800 19360 15940 19370
rect 15800 19320 15850 19360
rect 15890 19320 15940 19360
rect 15800 19310 15940 19320
rect 16020 19370 16050 19410
rect 16130 19370 16160 19410
rect 16020 19360 16160 19370
rect 16020 19320 16070 19360
rect 16110 19320 16160 19360
rect 16020 19310 16160 19320
rect 16240 19370 16270 19410
rect 16350 19370 16380 19410
rect 16240 19360 16380 19370
rect 16240 19320 16290 19360
rect 16330 19320 16380 19360
rect 16240 19310 16380 19320
rect 16460 19370 16490 19410
rect 16570 19370 16600 19410
rect 16460 19360 16600 19370
rect 16460 19320 16510 19360
rect 16550 19320 16600 19360
rect 16460 19310 16600 19320
rect 16680 19370 16710 19410
rect 16790 19370 16820 19410
rect 16680 19360 16820 19370
rect 16680 19320 16730 19360
rect 16770 19320 16820 19360
rect 16680 19310 16820 19320
rect 17090 19370 17120 19410
rect 17200 19370 17230 19410
rect 17090 19360 17230 19370
rect 17090 19320 17140 19360
rect 17180 19320 17230 19360
rect 17090 19310 17230 19320
rect 17310 19370 17340 19410
rect 17420 19370 17450 19410
rect 17310 19360 17450 19370
rect 17310 19320 17360 19360
rect 17400 19320 17450 19360
rect 17310 19310 17450 19320
rect 17530 19370 17560 19410
rect 17640 19370 17670 19410
rect 17530 19360 17670 19370
rect 17530 19320 17580 19360
rect 17620 19320 17670 19360
rect 17530 19310 17670 19320
rect 17750 19370 17780 19410
rect 17860 19370 17890 19410
rect 17750 19360 17890 19370
rect 17750 19320 17800 19360
rect 17840 19320 17890 19360
rect 17750 19310 17890 19320
rect 17970 19370 18000 19410
rect 18080 19370 18110 19410
rect 17970 19360 18110 19370
rect 17970 19320 18020 19360
rect 18060 19320 18110 19360
rect 17970 19310 18110 19320
rect 18190 19370 18220 19410
rect 18300 19370 18330 19410
rect 18190 19360 18330 19370
rect 18190 19320 18240 19360
rect 18280 19320 18330 19360
rect 18190 19310 18330 19320
rect 18410 19370 18440 19410
rect 18520 19370 18550 19410
rect 18410 19360 18550 19370
rect 18410 19320 18460 19360
rect 18500 19320 18550 19360
rect 18410 19310 18550 19320
rect 18630 19370 18660 19410
rect 18740 19370 18770 19410
rect 18630 19360 18770 19370
rect 18630 19320 18680 19360
rect 18720 19320 18770 19360
rect 18630 19310 18770 19320
rect 18850 19370 18880 19410
rect 18960 19370 18990 19410
rect 18850 19360 18990 19370
rect 18850 19320 18900 19360
rect 18940 19320 18990 19360
rect 18850 19310 18990 19320
rect 19070 19370 19100 19410
rect 19180 19370 19210 19410
rect 19070 19360 19210 19370
rect 19070 19320 19120 19360
rect 19160 19320 19210 19360
rect 19070 19310 19210 19320
rect 19290 19370 19320 19410
rect 19400 19370 19430 19410
rect 19290 19360 19430 19370
rect 19290 19320 19340 19360
rect 19380 19320 19430 19360
rect 19290 19310 19430 19320
rect 19510 19370 19540 19410
rect 19620 19370 19650 19410
rect 19510 19360 19650 19370
rect 19510 19320 19560 19360
rect 19600 19320 19650 19360
rect 19510 19310 19650 19320
rect 19730 19370 19760 19410
rect 19840 19370 19870 19410
rect 19730 19360 19870 19370
rect 19730 19320 19780 19360
rect 19820 19320 19870 19360
rect 19730 19310 19870 19320
rect 19950 19370 19980 19410
rect 20060 19370 20090 19410
rect 19950 19360 20090 19370
rect 19950 19320 20000 19360
rect 20040 19320 20090 19360
rect 19950 19310 20090 19320
rect 20170 19370 20200 19410
rect 20280 19370 20310 19410
rect 20170 19360 20310 19370
rect 20170 19320 20220 19360
rect 20260 19320 20310 19360
rect 20170 19310 20310 19320
rect 20390 19370 20420 19410
rect 20500 19370 20530 19410
rect 20390 19360 20530 19370
rect 20390 19320 20440 19360
rect 20480 19320 20530 19360
rect 20390 19310 20530 19320
rect 13740 19290 13880 19300
rect 14080 18470 14220 18480
rect 13180 18450 13320 18460
rect 13180 18410 13230 18450
rect 13270 18410 13320 18450
rect 13180 18400 13320 18410
rect 13180 18370 13210 18400
rect 12890 18350 12980 18370
rect 12890 18310 12900 18350
rect 12940 18310 12980 18350
rect 12890 18290 12980 18310
rect 13120 18350 13210 18370
rect 13120 18310 13130 18350
rect 13170 18330 13210 18350
rect 13290 18330 13320 18400
rect 13520 18450 13660 18460
rect 13520 18410 13570 18450
rect 13610 18410 13660 18450
rect 13520 18400 13660 18410
rect 13520 18370 13550 18400
rect 13170 18310 13320 18330
rect 13120 18290 13320 18310
rect 13460 18350 13550 18370
rect 13460 18310 13470 18350
rect 13510 18330 13550 18350
rect 13630 18330 13660 18400
rect 13740 18450 13880 18460
rect 13740 18410 13790 18450
rect 13830 18410 13880 18450
rect 13740 18400 13880 18410
rect 13740 18330 13770 18400
rect 13850 18330 13880 18400
rect 14080 18430 14130 18470
rect 14170 18430 14220 18470
rect 14080 18420 14220 18430
rect 14080 18370 14110 18420
rect 13510 18310 13880 18330
rect 13460 18290 13880 18310
rect 14020 18350 14110 18370
rect 14020 18310 14030 18350
rect 14070 18330 14110 18350
rect 14190 18330 14220 18420
rect 14300 18470 14440 18480
rect 14300 18430 14350 18470
rect 14390 18430 14440 18470
rect 14300 18420 14440 18430
rect 14300 18330 14330 18420
rect 14410 18330 14440 18420
rect 14520 18470 14660 18480
rect 14520 18430 14570 18470
rect 14610 18430 14660 18470
rect 14520 18420 14660 18430
rect 14520 18330 14550 18420
rect 14630 18330 14660 18420
rect 14740 18470 14880 18480
rect 14740 18430 14790 18470
rect 14830 18430 14880 18470
rect 14740 18420 14880 18430
rect 14740 18330 14770 18420
rect 14850 18330 14880 18420
rect 15140 18470 15280 18480
rect 15140 18430 15190 18470
rect 15230 18430 15280 18470
rect 15140 18420 15280 18430
rect 15140 18370 15170 18420
rect 14070 18310 14880 18330
rect 14020 18290 14880 18310
rect 15080 18350 15170 18370
rect 15080 18310 15090 18350
rect 15130 18330 15170 18350
rect 15250 18330 15280 18420
rect 15360 18470 15500 18480
rect 15360 18430 15410 18470
rect 15450 18430 15500 18470
rect 15360 18420 15500 18430
rect 15360 18330 15390 18420
rect 15470 18330 15500 18420
rect 15580 18470 15720 18480
rect 15580 18430 15630 18470
rect 15670 18430 15720 18470
rect 15580 18420 15720 18430
rect 15580 18330 15610 18420
rect 15690 18330 15720 18420
rect 15800 18470 15940 18480
rect 15800 18430 15850 18470
rect 15890 18430 15940 18470
rect 15800 18420 15940 18430
rect 15800 18330 15830 18420
rect 15910 18330 15940 18420
rect 16020 18470 16160 18480
rect 16020 18430 16070 18470
rect 16110 18430 16160 18470
rect 16020 18420 16160 18430
rect 16020 18330 16050 18420
rect 16130 18330 16160 18420
rect 16240 18470 16380 18480
rect 16240 18430 16290 18470
rect 16330 18430 16380 18470
rect 16240 18420 16380 18430
rect 16240 18330 16270 18420
rect 16350 18330 16380 18420
rect 16460 18470 16600 18480
rect 16460 18430 16510 18470
rect 16550 18430 16600 18470
rect 16460 18420 16600 18430
rect 16460 18330 16490 18420
rect 16570 18330 16600 18420
rect 16680 18470 16820 18480
rect 16680 18430 16730 18470
rect 16770 18430 16820 18470
rect 16680 18420 16820 18430
rect 16680 18330 16710 18420
rect 16790 18330 16820 18420
rect 17090 18470 17230 18480
rect 17090 18430 17140 18470
rect 17180 18430 17230 18470
rect 17090 18420 17230 18430
rect 17090 18370 17120 18420
rect 15130 18310 16820 18330
rect 15080 18290 16820 18310
rect 17020 18350 17120 18370
rect 17020 18310 17040 18350
rect 17080 18330 17120 18350
rect 17200 18330 17230 18420
rect 17310 18470 17450 18480
rect 17310 18430 17360 18470
rect 17400 18430 17450 18470
rect 17310 18420 17450 18430
rect 17310 18330 17340 18420
rect 17420 18330 17450 18420
rect 17530 18470 17670 18480
rect 17530 18430 17580 18470
rect 17620 18430 17670 18470
rect 17530 18420 17670 18430
rect 17530 18330 17560 18420
rect 17640 18330 17670 18420
rect 17750 18470 17890 18480
rect 17750 18430 17800 18470
rect 17840 18430 17890 18470
rect 17750 18420 17890 18430
rect 17750 18330 17780 18420
rect 17860 18330 17890 18420
rect 17970 18470 18110 18480
rect 17970 18430 18020 18470
rect 18060 18430 18110 18470
rect 17970 18420 18110 18430
rect 17970 18330 18000 18420
rect 18080 18330 18110 18420
rect 18190 18470 18330 18480
rect 18190 18430 18240 18470
rect 18280 18430 18330 18470
rect 18190 18420 18330 18430
rect 18190 18330 18220 18420
rect 18300 18330 18330 18420
rect 18410 18470 18550 18480
rect 18410 18430 18460 18470
rect 18500 18430 18550 18470
rect 18410 18420 18550 18430
rect 18410 18330 18440 18420
rect 18520 18330 18550 18420
rect 18630 18470 18770 18480
rect 18630 18430 18680 18470
rect 18720 18430 18770 18470
rect 18630 18420 18770 18430
rect 18630 18330 18660 18420
rect 18740 18330 18770 18420
rect 18850 18470 18990 18480
rect 18850 18430 18900 18470
rect 18940 18430 18990 18470
rect 18850 18420 18990 18430
rect 18850 18330 18880 18420
rect 18960 18330 18990 18420
rect 19070 18470 19210 18480
rect 19070 18430 19120 18470
rect 19160 18430 19210 18470
rect 19070 18420 19210 18430
rect 19070 18330 19100 18420
rect 19180 18330 19210 18420
rect 19290 18470 19430 18480
rect 19290 18430 19340 18470
rect 19380 18430 19430 18470
rect 19290 18420 19430 18430
rect 19290 18330 19320 18420
rect 19400 18330 19430 18420
rect 19510 18470 19650 18480
rect 19510 18430 19560 18470
rect 19600 18430 19650 18470
rect 19510 18420 19650 18430
rect 19510 18330 19540 18420
rect 19620 18330 19650 18420
rect 19730 18470 19870 18480
rect 19730 18430 19780 18470
rect 19820 18430 19870 18470
rect 19730 18420 19870 18430
rect 19730 18330 19760 18420
rect 19840 18330 19870 18420
rect 19950 18470 20090 18480
rect 19950 18430 20000 18470
rect 20040 18430 20090 18470
rect 19950 18420 20090 18430
rect 19950 18330 19980 18420
rect 20060 18330 20090 18420
rect 20170 18470 20310 18480
rect 20170 18430 20220 18470
rect 20260 18430 20310 18470
rect 20170 18420 20310 18430
rect 20170 18330 20200 18420
rect 20280 18330 20310 18420
rect 20390 18470 20530 18480
rect 20390 18430 20440 18470
rect 20480 18430 20530 18470
rect 20390 18420 20530 18430
rect 20390 18330 20420 18420
rect 20500 18330 20530 18420
rect 17080 18310 20530 18330
rect 17020 18290 20530 18310
rect 12950 18250 12980 18290
rect 13180 18250 13210 18290
rect 13290 18250 13320 18290
rect 13520 18250 13550 18290
rect 13630 18250 13660 18290
rect 13740 18250 13770 18290
rect 13850 18250 13880 18290
rect 14080 18250 14110 18290
rect 14190 18250 14220 18290
rect 14300 18250 14330 18290
rect 14410 18250 14440 18290
rect 14520 18250 14550 18290
rect 14630 18250 14660 18290
rect 14740 18250 14770 18290
rect 14850 18250 14880 18290
rect 15140 18250 15170 18290
rect 15250 18250 15280 18290
rect 15360 18250 15390 18290
rect 15470 18250 15500 18290
rect 15580 18250 15610 18290
rect 15690 18250 15720 18290
rect 15800 18250 15830 18290
rect 15910 18250 15940 18290
rect 16020 18250 16050 18290
rect 16130 18250 16160 18290
rect 16240 18250 16270 18290
rect 16350 18250 16380 18290
rect 16460 18250 16490 18290
rect 16570 18250 16600 18290
rect 16680 18250 16710 18290
rect 16790 18250 16820 18290
rect 17090 18250 17120 18290
rect 17200 18250 17230 18290
rect 17310 18250 17340 18290
rect 17420 18250 17450 18290
rect 17530 18250 17560 18290
rect 17640 18250 17670 18290
rect 17750 18250 17780 18290
rect 17860 18250 17890 18290
rect 17970 18250 18000 18290
rect 18080 18250 18110 18290
rect 18190 18250 18220 18290
rect 18300 18250 18330 18290
rect 18410 18250 18440 18290
rect 18520 18250 18550 18290
rect 18630 18250 18660 18290
rect 18740 18250 18770 18290
rect 18850 18250 18880 18290
rect 18960 18250 18990 18290
rect 19070 18250 19100 18290
rect 19180 18250 19210 18290
rect 19290 18250 19320 18290
rect 19400 18250 19430 18290
rect 19510 18250 19540 18290
rect 19620 18250 19650 18290
rect 19730 18250 19760 18290
rect 19840 18250 19870 18290
rect 19950 18250 19980 18290
rect 20060 18250 20090 18290
rect 20170 18250 20200 18290
rect 20280 18250 20310 18290
rect 20390 18250 20420 18290
rect 20500 18250 20530 18290
rect 12600 18220 12740 18250
rect 12600 17970 12630 18220
rect 12710 17970 12740 18220
rect 12950 18020 12980 18050
rect 13180 18020 13210 18050
rect 13290 18020 13320 18050
rect 13520 18020 13550 18050
rect 13630 18020 13660 18050
rect 13740 18020 13770 18050
rect 13850 18020 13880 18050
rect 14080 18020 14110 18050
rect 14190 18020 14220 18050
rect 14300 18020 14330 18050
rect 14410 18020 14440 18050
rect 14520 18020 14550 18050
rect 14630 18020 14660 18050
rect 14740 18020 14770 18050
rect 14850 18020 14880 18050
rect 15140 18020 15170 18050
rect 15250 18020 15280 18050
rect 15360 18020 15390 18050
rect 15470 18020 15500 18050
rect 15580 18020 15610 18050
rect 15690 18020 15720 18050
rect 15800 18020 15830 18050
rect 15910 18020 15940 18050
rect 16020 18020 16050 18050
rect 16130 18020 16160 18050
rect 16240 18020 16270 18050
rect 16350 18020 16380 18050
rect 16460 18020 16490 18050
rect 16570 18020 16600 18050
rect 16680 18020 16710 18050
rect 16790 18020 16820 18050
rect 17090 18020 17120 18050
rect 17200 18020 17230 18050
rect 17310 18020 17340 18050
rect 17420 18020 17450 18050
rect 17530 18020 17560 18050
rect 17640 18020 17670 18050
rect 17750 18020 17780 18050
rect 17860 18020 17890 18050
rect 17970 18020 18000 18050
rect 18080 18020 18110 18050
rect 18190 18020 18220 18050
rect 18300 18020 18330 18050
rect 18410 18020 18440 18050
rect 18520 18020 18550 18050
rect 18630 18020 18660 18050
rect 18740 18020 18770 18050
rect 18850 18020 18880 18050
rect 18960 18020 18990 18050
rect 19070 18020 19100 18050
rect 19180 18020 19210 18050
rect 19290 18020 19320 18050
rect 19400 18020 19430 18050
rect 19510 18020 19540 18050
rect 19620 18020 19650 18050
rect 19730 18020 19760 18050
rect 19840 18020 19870 18050
rect 19950 18020 19980 18050
rect 20060 18020 20090 18050
rect 20170 18020 20200 18050
rect 20280 18020 20310 18050
rect 20390 18020 20420 18050
rect 20500 18020 20530 18050
rect 8550 17740 8580 17770
rect 8700 17740 8730 17770
rect 9290 17740 9320 17770
rect 9400 17740 9430 17770
rect 9630 17740 9660 17770
rect 9740 17740 9770 17770
rect 9890 17740 9920 17770
rect 10000 17740 10030 17770
rect 10230 17740 10260 17770
rect 10340 17740 10370 17770
rect 10620 17740 10650 17770
rect 10730 17740 10760 17770
rect 10880 17740 10910 17770
rect 10990 17740 11020 17770
rect 11220 17740 11250 17770
rect 11330 17740 11360 17770
rect 11620 17740 11650 17770
rect 11730 17740 11760 17770
rect 11880 17740 11910 17770
rect 11990 17740 12020 17770
rect 12220 17740 12250 17770
rect 12330 17740 12360 17770
rect 12600 17740 12630 17770
rect 12710 17740 12740 17770
rect 9830 15550 9860 15580
rect 9940 15550 9970 15580
rect 10370 15550 10400 15580
rect 10480 15550 10510 15580
rect 10630 15550 10660 15580
rect 10740 15550 10770 15580
rect 10970 15550 11000 15580
rect 11080 15550 11110 15580
rect 11360 15550 11390 15580
rect 11470 15550 11500 15580
rect 11620 15550 11650 15580
rect 11730 15550 11760 15580
rect 11960 15550 11990 15580
rect 12070 15550 12100 15580
rect 12360 15550 12390 15580
rect 12470 15550 12500 15580
rect 12620 15550 12650 15580
rect 12730 15550 12760 15580
rect 12960 15550 12990 15580
rect 13070 15550 13100 15580
rect 9830 15330 9860 15350
rect 9940 15330 9970 15350
rect 9830 15300 9970 15330
rect 9830 15120 9860 15300
rect 9730 15110 9860 15120
rect 9730 15050 9750 15110
rect 9810 15050 9860 15110
rect 9730 15040 9860 15050
rect 9830 14910 9860 15040
rect 9940 15010 9970 15300
rect 10370 15030 10400 15150
rect 10260 15020 10400 15030
rect 10260 14960 10280 15020
rect 10350 15000 10400 15020
rect 10480 15000 10510 15150
rect 10630 15130 10660 15150
rect 10570 15110 10660 15130
rect 10570 15070 10580 15110
rect 10620 15100 10660 15110
rect 10740 15100 10770 15150
rect 10620 15070 10770 15100
rect 10570 15050 10660 15070
rect 10350 14970 10510 15000
rect 10350 14960 10400 14970
rect 10260 14950 10400 14960
rect 9940 14910 9970 14950
rect 10370 14910 10400 14950
rect 10480 14910 10510 14970
rect 10630 14910 10660 15050
rect 10740 14910 10770 15070
rect 10970 15010 11000 15350
rect 11080 15010 11110 15350
rect 11360 15030 11390 15150
rect 11300 15010 11390 15030
rect 10880 15000 11000 15010
rect 10880 14960 10900 15000
rect 10940 14960 11000 15000
rect 10880 14950 11000 14960
rect 11300 14970 11310 15010
rect 11350 15000 11390 15010
rect 11470 15000 11500 15150
rect 11620 15130 11650 15150
rect 11560 15110 11650 15130
rect 11560 15070 11570 15110
rect 11610 15100 11650 15110
rect 11730 15100 11760 15150
rect 11610 15070 11760 15100
rect 11560 15050 11650 15070
rect 11350 14970 11500 15000
rect 11300 14950 11390 14970
rect 10970 14910 11000 14950
rect 11080 14910 11110 14950
rect 11360 14910 11390 14950
rect 11470 14910 11500 14970
rect 11620 14910 11650 15050
rect 11730 14910 11760 15070
rect 11960 15010 11990 15350
rect 12070 15010 12100 15350
rect 12360 15030 12390 15150
rect 12300 15010 12390 15030
rect 11870 15000 11990 15010
rect 11870 14960 11890 15000
rect 11930 14960 11990 15000
rect 11870 14950 11990 14960
rect 12300 14970 12310 15010
rect 12350 15000 12390 15010
rect 12470 15000 12500 15150
rect 12620 15130 12650 15150
rect 12560 15110 12650 15130
rect 12560 15070 12570 15110
rect 12610 15100 12650 15110
rect 12730 15100 12760 15150
rect 12610 15070 12760 15100
rect 12560 15050 12650 15070
rect 12350 14970 12500 15000
rect 12300 14950 12390 14970
rect 11960 14910 11990 14950
rect 12070 14910 12100 14950
rect 12360 14910 12390 14950
rect 12470 14910 12500 14970
rect 12620 14910 12650 15050
rect 12730 14910 12760 15070
rect 12960 15010 12990 15350
rect 13070 15010 13100 15350
rect 13310 15270 13340 15300
rect 13540 15270 13570 15300
rect 13650 15270 13680 15300
rect 13880 15270 13910 15300
rect 13990 15270 14020 15300
rect 14100 15270 14130 15300
rect 14210 15270 14240 15300
rect 14440 15270 14470 15300
rect 14550 15270 14580 15300
rect 14660 15270 14690 15300
rect 14770 15270 14800 15300
rect 14880 15270 14910 15300
rect 14990 15270 15020 15300
rect 15100 15270 15130 15300
rect 15210 15270 15240 15300
rect 15500 15270 15530 15300
rect 15610 15270 15640 15300
rect 15720 15270 15750 15300
rect 15830 15270 15860 15300
rect 15940 15270 15970 15300
rect 16050 15270 16080 15300
rect 16160 15270 16190 15300
rect 16270 15270 16300 15300
rect 16380 15270 16410 15300
rect 16490 15270 16520 15300
rect 16600 15270 16630 15300
rect 16710 15270 16740 15300
rect 16820 15270 16850 15300
rect 16930 15270 16960 15300
rect 17040 15270 17070 15300
rect 17150 15270 17180 15300
rect 17450 15270 17480 15300
rect 17560 15270 17590 15300
rect 17670 15270 17700 15300
rect 17780 15270 17810 15300
rect 17890 15270 17920 15300
rect 18000 15270 18030 15300
rect 18110 15270 18140 15300
rect 18220 15270 18250 15300
rect 18330 15270 18360 15300
rect 18440 15270 18470 15300
rect 18550 15270 18580 15300
rect 18660 15270 18690 15300
rect 18770 15270 18800 15300
rect 18880 15270 18910 15300
rect 18990 15270 19020 15300
rect 19100 15270 19130 15300
rect 19210 15270 19240 15300
rect 19320 15270 19350 15300
rect 19430 15270 19460 15300
rect 19540 15270 19570 15300
rect 19650 15270 19680 15300
rect 19760 15270 19790 15300
rect 19870 15270 19900 15300
rect 19980 15270 20010 15300
rect 20090 15270 20120 15300
rect 20200 15270 20230 15300
rect 20310 15270 20340 15300
rect 20420 15270 20450 15300
rect 20530 15270 20560 15300
rect 20640 15270 20670 15300
rect 20750 15270 20780 15300
rect 20860 15270 20890 15300
rect 13310 15030 13340 15070
rect 13540 15030 13570 15070
rect 13650 15030 13680 15070
rect 13880 15030 13910 15070
rect 13990 15030 14020 15070
rect 14100 15030 14130 15070
rect 14210 15030 14240 15070
rect 14440 15030 14470 15070
rect 14550 15030 14580 15070
rect 14660 15030 14690 15070
rect 14770 15030 14800 15070
rect 14880 15030 14910 15070
rect 14990 15030 15020 15070
rect 15100 15030 15130 15070
rect 15210 15030 15240 15070
rect 15500 15030 15530 15070
rect 15610 15030 15640 15070
rect 15720 15030 15750 15070
rect 15830 15030 15860 15070
rect 15940 15030 15970 15070
rect 16050 15030 16080 15070
rect 16160 15030 16190 15070
rect 16270 15030 16300 15070
rect 16380 15030 16410 15070
rect 16490 15030 16520 15070
rect 16600 15030 16630 15070
rect 16710 15030 16740 15070
rect 16820 15030 16850 15070
rect 16930 15030 16960 15070
rect 17040 15030 17070 15070
rect 17150 15030 17180 15070
rect 17450 15030 17480 15070
rect 17560 15030 17590 15070
rect 17670 15030 17700 15070
rect 17780 15030 17810 15070
rect 17890 15030 17920 15070
rect 18000 15030 18030 15070
rect 18110 15030 18140 15070
rect 18220 15030 18250 15070
rect 18330 15030 18360 15070
rect 18440 15030 18470 15070
rect 18550 15030 18580 15070
rect 18660 15030 18690 15070
rect 18770 15030 18800 15070
rect 18880 15030 18910 15070
rect 18990 15030 19020 15070
rect 19100 15030 19130 15070
rect 19210 15030 19240 15070
rect 19320 15030 19350 15070
rect 19430 15030 19460 15070
rect 19540 15030 19570 15070
rect 19650 15030 19680 15070
rect 19760 15030 19790 15070
rect 19870 15030 19900 15070
rect 19980 15030 20010 15070
rect 20090 15030 20120 15070
rect 20200 15030 20230 15070
rect 20310 15030 20340 15070
rect 20420 15030 20450 15070
rect 20530 15030 20560 15070
rect 20640 15030 20670 15070
rect 20750 15030 20780 15070
rect 20860 15030 20890 15070
rect 13250 15010 13340 15030
rect 12870 15000 12990 15010
rect 12870 14960 12890 15000
rect 12930 14960 12990 15000
rect 12870 14950 12990 14960
rect 13250 14970 13260 15010
rect 13300 14970 13340 15010
rect 13250 14950 13340 14970
rect 13480 15010 13680 15030
rect 13480 14970 13490 15010
rect 13530 14990 13680 15010
rect 13530 14970 13570 14990
rect 13480 14950 13570 14970
rect 12960 14910 12990 14950
rect 13070 14910 13100 14950
rect 13310 14910 13340 14950
rect 13540 14910 13570 14950
rect 13650 14910 13680 14990
rect 13820 15010 14240 15030
rect 13820 14970 13830 15010
rect 13870 14990 14240 15010
rect 13870 14970 13910 14990
rect 13820 14950 13910 14970
rect 13880 14910 13910 14950
rect 13990 14910 14020 14990
rect 14100 14910 14130 14990
rect 14210 14910 14240 14990
rect 14380 15010 15240 15030
rect 14380 14970 14390 15010
rect 14430 14990 15240 15010
rect 14430 14970 14470 14990
rect 14380 14950 14470 14970
rect 14440 14910 14470 14950
rect 14550 14910 14580 14990
rect 14660 14910 14690 14990
rect 14770 14910 14800 14990
rect 14880 14910 14910 14990
rect 14990 14910 15020 14990
rect 15100 14910 15130 14990
rect 15210 14910 15240 14990
rect 15440 15010 17180 15030
rect 15440 14970 15450 15010
rect 15490 14990 17180 15010
rect 15490 14970 15530 14990
rect 15440 14950 15530 14970
rect 15500 14910 15530 14950
rect 15610 14910 15640 14990
rect 15720 14910 15750 14990
rect 15830 14910 15860 14990
rect 15940 14910 15970 14990
rect 16050 14910 16080 14990
rect 16160 14910 16190 14990
rect 16270 14910 16300 14990
rect 16380 14910 16410 14990
rect 16490 14910 16520 14990
rect 16600 14910 16630 14990
rect 16710 14910 16740 14990
rect 16820 14910 16850 14990
rect 16930 14910 16960 14990
rect 17040 14910 17070 14990
rect 17150 14910 17180 14990
rect 17380 15010 20890 15030
rect 17380 14970 17400 15010
rect 17440 14990 20890 15010
rect 17440 14970 17480 14990
rect 17380 14950 17480 14970
rect 17450 14910 17480 14950
rect 17560 14910 17590 14990
rect 17670 14910 17700 14990
rect 17780 14910 17810 14990
rect 17890 14910 17920 14990
rect 18000 14910 18030 14990
rect 18110 14910 18140 14990
rect 18220 14910 18250 14990
rect 18330 14910 18360 14990
rect 18440 14910 18470 14990
rect 18550 14910 18580 14990
rect 18660 14910 18690 14990
rect 18770 14910 18800 14990
rect 18880 14910 18910 14990
rect 18990 14910 19020 14990
rect 19100 14910 19130 14990
rect 19210 14910 19240 14990
rect 19320 14910 19350 14990
rect 19430 14910 19460 14990
rect 19540 14910 19570 14990
rect 19650 14910 19680 14990
rect 19760 14910 19790 14990
rect 19870 14910 19900 14990
rect 19980 14910 20010 14990
rect 20090 14910 20120 14990
rect 20200 14910 20230 14990
rect 20310 14910 20340 14990
rect 20420 14910 20450 14990
rect 20530 14910 20560 14990
rect 20640 14910 20670 14990
rect 20750 14910 20780 14990
rect 20860 14910 20890 14990
rect 9830 14380 9860 14410
rect 9940 14380 9970 14410
rect 10370 14380 10400 14410
rect 10480 14380 10510 14410
rect 10630 14380 10660 14410
rect 10740 14380 10770 14410
rect 10970 14380 11000 14410
rect 11080 14380 11110 14410
rect 11360 14380 11390 14410
rect 11470 14380 11500 14410
rect 11620 14380 11650 14410
rect 11730 14380 11760 14410
rect 11960 14380 11990 14410
rect 12070 14380 12100 14410
rect 12360 14380 12390 14410
rect 12470 14380 12500 14410
rect 12620 14380 12650 14410
rect 12730 14380 12760 14410
rect 12960 14380 12990 14410
rect 13070 14380 13100 14410
rect 13310 14380 13340 14410
rect 13540 14380 13570 14410
rect 13650 14380 13680 14410
rect 13880 14380 13910 14410
rect 13990 14380 14020 14410
rect 14100 14380 14130 14410
rect 14210 14380 14240 14410
rect 14440 14380 14470 14410
rect 14550 14380 14580 14410
rect 14660 14380 14690 14410
rect 14770 14380 14800 14410
rect 14880 14380 14910 14410
rect 14990 14380 15020 14410
rect 15100 14380 15130 14410
rect 15210 14380 15240 14410
rect 15500 14380 15530 14410
rect 15610 14380 15640 14410
rect 15720 14380 15750 14410
rect 15830 14380 15860 14410
rect 15940 14380 15970 14410
rect 16050 14380 16080 14410
rect 16160 14380 16190 14410
rect 16270 14380 16300 14410
rect 16380 14380 16410 14410
rect 16490 14380 16520 14410
rect 16600 14380 16630 14410
rect 16710 14380 16740 14410
rect 16820 14380 16850 14410
rect 16930 14380 16960 14410
rect 17040 14380 17070 14410
rect 17150 14380 17180 14410
rect 17450 14380 17480 14410
rect 17560 14380 17590 14410
rect 17670 14380 17700 14410
rect 17780 14380 17810 14410
rect 17890 14380 17920 14410
rect 18000 14380 18030 14410
rect 18110 14380 18140 14410
rect 18220 14380 18250 14410
rect 18330 14380 18360 14410
rect 18440 14380 18470 14410
rect 18550 14380 18580 14410
rect 18660 14380 18690 14410
rect 18770 14380 18800 14410
rect 18880 14380 18910 14410
rect 18990 14380 19020 14410
rect 19100 14380 19130 14410
rect 19210 14380 19240 14410
rect 19320 14380 19350 14410
rect 19430 14380 19460 14410
rect 19540 14380 19570 14410
rect 19650 14380 19680 14410
rect 19760 14380 19790 14410
rect 19870 14380 19900 14410
rect 19980 14380 20010 14410
rect 20090 14380 20120 14410
rect 20200 14380 20230 14410
rect 20310 14380 20340 14410
rect 20420 14380 20450 14410
rect 20530 14380 20560 14410
rect 20640 14380 20670 14410
rect 20750 14380 20780 14410
rect 20860 14380 20890 14410
rect 7350 13260 7380 13290
rect 7460 13260 7490 13290
rect 7870 13260 7900 13290
rect 7980 13260 8010 13290
rect 8130 13260 8160 13290
rect 8240 13260 8270 13290
rect 8620 13260 8650 13290
rect 8770 13260 8800 13290
rect 9000 13260 9030 13290
rect 9260 13260 9290 13290
rect 9510 13260 9540 13290
rect 9930 13260 9960 13290
rect 10040 13260 10070 13290
rect 10470 13260 10500 13290
rect 10580 13260 10610 13290
rect 10730 13260 10760 13290
rect 10840 13260 10870 13290
rect 11070 13260 11100 13290
rect 11180 13260 11210 13290
rect 11460 13260 11490 13290
rect 11570 13260 11600 13290
rect 11720 13260 11750 13290
rect 11830 13260 11860 13290
rect 12060 13260 12090 13290
rect 12170 13260 12200 13290
rect 12460 13260 12490 13290
rect 12570 13260 12600 13290
rect 12720 13260 12750 13290
rect 12830 13260 12860 13290
rect 13060 13260 13090 13290
rect 13170 13260 13200 13290
rect 13410 13260 13440 13290
rect 13640 13260 13670 13290
rect 13750 13260 13780 13290
rect 13980 13260 14010 13290
rect 14090 13260 14120 13290
rect 14200 13260 14230 13290
rect 14310 13260 14340 13290
rect 14540 13260 14570 13290
rect 14650 13260 14680 13290
rect 14760 13260 14790 13290
rect 14870 13260 14900 13290
rect 14980 13260 15010 13290
rect 15090 13260 15120 13290
rect 15200 13260 15230 13290
rect 15310 13260 15340 13290
rect 15600 13260 15630 13290
rect 15710 13260 15740 13290
rect 15820 13260 15850 13290
rect 15930 13260 15960 13290
rect 16040 13260 16070 13290
rect 16150 13260 16180 13290
rect 16260 13260 16290 13290
rect 16370 13260 16400 13290
rect 16480 13260 16510 13290
rect 16590 13260 16620 13290
rect 16700 13260 16730 13290
rect 16810 13260 16840 13290
rect 16920 13260 16950 13290
rect 17030 13260 17060 13290
rect 17140 13260 17170 13290
rect 17250 13260 17280 13290
rect 17550 13260 17580 13290
rect 17660 13260 17690 13290
rect 17770 13260 17800 13290
rect 17880 13260 17910 13290
rect 17990 13260 18020 13290
rect 18100 13260 18130 13290
rect 18210 13260 18240 13290
rect 18320 13260 18350 13290
rect 18430 13260 18460 13290
rect 18540 13260 18570 13290
rect 18650 13260 18680 13290
rect 18760 13260 18790 13290
rect 18870 13260 18900 13290
rect 18980 13260 19010 13290
rect 19090 13260 19120 13290
rect 19200 13260 19230 13290
rect 19310 13260 19340 13290
rect 19420 13260 19450 13290
rect 19530 13260 19560 13290
rect 19640 13260 19670 13290
rect 19750 13260 19780 13290
rect 19860 13260 19890 13290
rect 19970 13260 20000 13290
rect 20080 13260 20110 13290
rect 20190 13260 20220 13290
rect 20300 13260 20330 13290
rect 20410 13260 20440 13290
rect 20520 13260 20550 13290
rect 20630 13260 20660 13290
rect 20740 13260 20770 13290
rect 20850 13260 20880 13290
rect 20960 13260 20990 13290
rect 7350 12720 7380 12760
rect 7250 12710 7380 12720
rect 7250 12650 7270 12710
rect 7330 12650 7380 12710
rect 7250 12640 7380 12650
rect 7350 12380 7380 12640
rect 7460 12380 7490 12760
rect 7870 12720 7900 12760
rect 7800 12700 7900 12720
rect 7980 12700 8010 12760
rect 7800 12660 7820 12700
rect 7860 12670 8010 12700
rect 7860 12660 7900 12670
rect 7800 12640 7900 12660
rect 7870 12520 7900 12640
rect 7980 12520 8010 12670
rect 8130 12620 8160 12760
rect 8070 12600 8160 12620
rect 8240 12600 8270 12760
rect 8620 12710 8650 12760
rect 8550 12690 8650 12710
rect 8550 12650 8570 12690
rect 8610 12650 8650 12690
rect 8550 12630 8650 12650
rect 8070 12560 8080 12600
rect 8120 12570 8270 12600
rect 8120 12560 8160 12570
rect 8070 12540 8160 12560
rect 8130 12520 8160 12540
rect 8240 12520 8270 12570
rect 7350 12350 7490 12380
rect 7350 12320 7380 12350
rect 7460 12320 7490 12350
rect 8620 12480 8650 12630
rect 8770 12600 8800 12760
rect 9000 12720 9030 12760
rect 9260 12720 9290 12760
rect 9510 12720 9540 12760
rect 9930 12720 9960 12760
rect 10040 12720 10070 12760
rect 10470 12720 10500 12760
rect 8930 12700 9030 12720
rect 8930 12660 8950 12700
rect 8990 12660 9030 12700
rect 8930 12640 9030 12660
rect 9190 12700 9290 12720
rect 9190 12660 9210 12700
rect 9250 12660 9290 12700
rect 9190 12640 9290 12660
rect 9440 12700 9540 12720
rect 9440 12660 9460 12700
rect 9500 12660 9540 12700
rect 9840 12710 9960 12720
rect 9840 12670 9860 12710
rect 9900 12670 9960 12710
rect 9840 12660 9960 12670
rect 10410 12700 10500 12720
rect 10580 12700 10610 12760
rect 10410 12660 10420 12700
rect 10460 12670 10610 12700
rect 10460 12660 10500 12670
rect 9440 12640 9540 12660
rect 8700 12580 8800 12600
rect 9000 12590 9030 12640
rect 9260 12590 9290 12640
rect 9510 12590 9540 12640
rect 8700 12540 8720 12580
rect 8760 12540 8800 12580
rect 8700 12520 8800 12540
rect 8770 12480 8800 12520
rect 7350 12090 7380 12120
rect 7460 12090 7490 12120
rect 7870 12090 7900 12120
rect 7980 12090 8010 12120
rect 8130 12090 8160 12120
rect 8240 12090 8270 12120
rect 9000 12360 9030 12390
rect 9260 12360 9290 12390
rect 9510 12360 9540 12390
rect 9930 12370 9960 12660
rect 10040 12370 10070 12660
rect 10410 12640 10500 12660
rect 10470 12520 10500 12640
rect 10580 12520 10610 12670
rect 10730 12620 10760 12760
rect 10670 12600 10760 12620
rect 10840 12600 10870 12760
rect 11070 12720 11100 12760
rect 11180 12720 11210 12760
rect 11460 12720 11490 12760
rect 10980 12710 11100 12720
rect 10980 12670 11000 12710
rect 11040 12670 11100 12710
rect 10980 12660 11100 12670
rect 11400 12700 11490 12720
rect 11570 12700 11600 12760
rect 11400 12660 11410 12700
rect 11450 12670 11600 12700
rect 11450 12660 11490 12670
rect 10670 12560 10680 12600
rect 10720 12570 10870 12600
rect 10720 12560 10760 12570
rect 10670 12540 10760 12560
rect 10730 12520 10760 12540
rect 10840 12520 10870 12570
rect 9930 12340 10070 12370
rect 9930 12320 9960 12340
rect 10040 12320 10070 12340
rect 11070 12320 11100 12660
rect 11180 12320 11210 12660
rect 11400 12640 11490 12660
rect 11460 12520 11490 12640
rect 11570 12520 11600 12670
rect 11720 12620 11750 12760
rect 11660 12600 11750 12620
rect 11830 12600 11860 12760
rect 12060 12720 12090 12760
rect 12170 12720 12200 12760
rect 12460 12720 12490 12760
rect 11970 12710 12090 12720
rect 11970 12670 11990 12710
rect 12030 12670 12090 12710
rect 11970 12660 12090 12670
rect 12400 12700 12490 12720
rect 12570 12700 12600 12760
rect 12400 12660 12410 12700
rect 12450 12670 12600 12700
rect 12450 12660 12490 12670
rect 11660 12560 11670 12600
rect 11710 12570 11860 12600
rect 11710 12560 11750 12570
rect 11660 12540 11750 12560
rect 11720 12520 11750 12540
rect 11830 12520 11860 12570
rect 12060 12320 12090 12660
rect 12170 12320 12200 12660
rect 12400 12640 12490 12660
rect 12460 12520 12490 12640
rect 12570 12520 12600 12670
rect 12720 12620 12750 12760
rect 12660 12600 12750 12620
rect 12830 12600 12860 12760
rect 13060 12720 13090 12760
rect 13170 12720 13200 12760
rect 13410 12720 13440 12760
rect 13640 12720 13670 12760
rect 12970 12710 13090 12720
rect 12970 12670 12990 12710
rect 13030 12670 13090 12710
rect 12970 12660 13090 12670
rect 13350 12700 13440 12720
rect 13350 12660 13360 12700
rect 13400 12660 13440 12700
rect 12660 12560 12670 12600
rect 12710 12570 12860 12600
rect 12710 12560 12750 12570
rect 12660 12540 12750 12560
rect 12720 12520 12750 12540
rect 12830 12520 12860 12570
rect 13060 12320 13090 12660
rect 13170 12320 13200 12660
rect 13350 12640 13440 12660
rect 13580 12700 13670 12720
rect 13580 12660 13590 12700
rect 13630 12680 13670 12700
rect 13750 12680 13780 12760
rect 13980 12720 14010 12760
rect 13630 12660 13780 12680
rect 13580 12640 13780 12660
rect 13920 12700 14010 12720
rect 13920 12660 13930 12700
rect 13970 12680 14010 12700
rect 14090 12680 14120 12760
rect 14200 12680 14230 12760
rect 14310 12680 14340 12760
rect 14540 12720 14570 12760
rect 13970 12660 14340 12680
rect 13920 12640 14340 12660
rect 14480 12700 14570 12720
rect 14480 12660 14490 12700
rect 14530 12680 14570 12700
rect 14650 12680 14680 12760
rect 14760 12680 14790 12760
rect 14870 12680 14900 12760
rect 14980 12680 15010 12760
rect 15090 12680 15120 12760
rect 15200 12680 15230 12760
rect 15310 12680 15340 12760
rect 15600 12720 15630 12760
rect 14530 12660 15340 12680
rect 14480 12640 15340 12660
rect 15540 12700 15630 12720
rect 15540 12660 15550 12700
rect 15590 12680 15630 12700
rect 15710 12680 15740 12760
rect 15820 12680 15850 12760
rect 15930 12680 15960 12760
rect 16040 12680 16070 12760
rect 16150 12680 16180 12760
rect 16260 12680 16290 12760
rect 16370 12680 16400 12760
rect 16480 12680 16510 12760
rect 16590 12680 16620 12760
rect 16700 12680 16730 12760
rect 16810 12680 16840 12760
rect 16920 12680 16950 12760
rect 17030 12680 17060 12760
rect 17140 12680 17170 12760
rect 17250 12680 17280 12760
rect 17550 12720 17580 12760
rect 15590 12660 17280 12680
rect 15540 12640 17280 12660
rect 17480 12700 17580 12720
rect 17480 12660 17500 12700
rect 17540 12680 17580 12700
rect 17660 12680 17690 12760
rect 17770 12680 17800 12760
rect 17880 12680 17910 12760
rect 17990 12680 18020 12760
rect 18100 12680 18130 12760
rect 18210 12680 18240 12760
rect 18320 12680 18350 12760
rect 18430 12680 18460 12760
rect 18540 12680 18570 12760
rect 18650 12680 18680 12760
rect 18760 12680 18790 12760
rect 18870 12680 18900 12760
rect 18980 12680 19010 12760
rect 19090 12680 19120 12760
rect 19200 12680 19230 12760
rect 19310 12680 19340 12760
rect 19420 12680 19450 12760
rect 19530 12680 19560 12760
rect 19640 12680 19670 12760
rect 19750 12680 19780 12760
rect 19860 12680 19890 12760
rect 19970 12680 20000 12760
rect 20080 12680 20110 12760
rect 20190 12680 20220 12760
rect 20300 12680 20330 12760
rect 20410 12680 20440 12760
rect 20520 12680 20550 12760
rect 20630 12680 20660 12760
rect 20740 12680 20770 12760
rect 20850 12680 20880 12760
rect 20960 12680 20990 12760
rect 17540 12660 20990 12680
rect 17480 12640 20990 12660
rect 13410 12600 13440 12640
rect 13640 12600 13670 12640
rect 13750 12600 13780 12640
rect 13980 12600 14010 12640
rect 14090 12600 14120 12640
rect 14200 12600 14230 12640
rect 14310 12600 14340 12640
rect 14540 12600 14570 12640
rect 14650 12600 14680 12640
rect 14760 12600 14790 12640
rect 14870 12600 14900 12640
rect 14980 12600 15010 12640
rect 15090 12600 15120 12640
rect 15200 12600 15230 12640
rect 15310 12600 15340 12640
rect 15600 12600 15630 12640
rect 15710 12600 15740 12640
rect 15820 12600 15850 12640
rect 15930 12600 15960 12640
rect 16040 12600 16070 12640
rect 16150 12600 16180 12640
rect 16260 12600 16290 12640
rect 16370 12600 16400 12640
rect 16480 12600 16510 12640
rect 16590 12600 16620 12640
rect 16700 12600 16730 12640
rect 16810 12600 16840 12640
rect 16920 12600 16950 12640
rect 17030 12600 17060 12640
rect 17140 12600 17170 12640
rect 17250 12600 17280 12640
rect 17550 12600 17580 12640
rect 17660 12600 17690 12640
rect 17770 12600 17800 12640
rect 17880 12600 17910 12640
rect 17990 12600 18020 12640
rect 18100 12600 18130 12640
rect 18210 12600 18240 12640
rect 18320 12600 18350 12640
rect 18430 12600 18460 12640
rect 18540 12600 18570 12640
rect 18650 12600 18680 12640
rect 18760 12600 18790 12640
rect 18870 12600 18900 12640
rect 18980 12600 19010 12640
rect 19090 12600 19120 12640
rect 19200 12600 19230 12640
rect 19310 12600 19340 12640
rect 19420 12600 19450 12640
rect 19530 12600 19560 12640
rect 19640 12600 19670 12640
rect 19750 12600 19780 12640
rect 19860 12600 19890 12640
rect 19970 12600 20000 12640
rect 20080 12600 20110 12640
rect 20190 12600 20220 12640
rect 20300 12600 20330 12640
rect 20410 12600 20440 12640
rect 20520 12600 20550 12640
rect 20630 12600 20660 12640
rect 20740 12600 20770 12640
rect 20850 12600 20880 12640
rect 20960 12600 20990 12640
rect 13410 12370 13440 12400
rect 13640 12370 13670 12400
rect 13750 12370 13780 12400
rect 13980 12370 14010 12400
rect 14090 12370 14120 12400
rect 14200 12370 14230 12400
rect 14310 12370 14340 12400
rect 14540 12370 14570 12400
rect 14650 12370 14680 12400
rect 14760 12370 14790 12400
rect 14870 12370 14900 12400
rect 14980 12370 15010 12400
rect 15090 12370 15120 12400
rect 15200 12370 15230 12400
rect 15310 12370 15340 12400
rect 15600 12370 15630 12400
rect 15710 12370 15740 12400
rect 15820 12370 15850 12400
rect 15930 12370 15960 12400
rect 16040 12370 16070 12400
rect 16150 12370 16180 12400
rect 16260 12370 16290 12400
rect 16370 12370 16400 12400
rect 16480 12370 16510 12400
rect 16590 12370 16620 12400
rect 16700 12370 16730 12400
rect 16810 12370 16840 12400
rect 16920 12370 16950 12400
rect 17030 12370 17060 12400
rect 17140 12370 17170 12400
rect 17250 12370 17280 12400
rect 17550 12370 17580 12400
rect 17660 12370 17690 12400
rect 17770 12370 17800 12400
rect 17880 12370 17910 12400
rect 17990 12370 18020 12400
rect 18100 12370 18130 12400
rect 18210 12370 18240 12400
rect 18320 12370 18350 12400
rect 18430 12370 18460 12400
rect 18540 12370 18570 12400
rect 18650 12370 18680 12400
rect 18760 12370 18790 12400
rect 18870 12370 18900 12400
rect 18980 12370 19010 12400
rect 19090 12370 19120 12400
rect 19200 12370 19230 12400
rect 19310 12370 19340 12400
rect 19420 12370 19450 12400
rect 19530 12370 19560 12400
rect 19640 12370 19670 12400
rect 19750 12370 19780 12400
rect 19860 12370 19890 12400
rect 19970 12370 20000 12400
rect 20080 12370 20110 12400
rect 20190 12370 20220 12400
rect 20300 12370 20330 12400
rect 20410 12370 20440 12400
rect 20520 12370 20550 12400
rect 20630 12370 20660 12400
rect 20740 12370 20770 12400
rect 20850 12370 20880 12400
rect 20960 12370 20990 12400
rect 9930 12090 9960 12120
rect 10040 12090 10070 12120
rect 10470 12090 10500 12120
rect 10580 12090 10610 12120
rect 10730 12090 10760 12120
rect 10840 12090 10870 12120
rect 11070 12090 11100 12120
rect 11180 12090 11210 12120
rect 11460 12090 11490 12120
rect 11570 12090 11600 12120
rect 11720 12090 11750 12120
rect 11830 12090 11860 12120
rect 12060 12090 12090 12120
rect 12170 12090 12200 12120
rect 12460 12090 12490 12120
rect 12570 12090 12600 12120
rect 12720 12090 12750 12120
rect 12830 12090 12860 12120
rect 13060 12090 13090 12120
rect 13170 12090 13200 12120
rect 8620 12050 8650 12080
rect 8770 12050 8800 12080
rect 7920 11300 7950 11340
rect 8030 11300 8060 11340
rect 8180 11300 8210 11340
rect 8290 11300 8320 11340
rect 7350 10930 7380 10960
rect 7460 10930 7490 10960
rect 7920 10870 7950 11100
rect 7840 10850 7950 10870
rect 7840 10790 7850 10850
rect 7910 10840 7950 10850
rect 8030 10840 8060 11100
rect 8180 10960 8210 11100
rect 8120 10940 8210 10960
rect 8290 10940 8320 11100
rect 8710 10980 8740 11010
rect 8860 10980 8890 11010
rect 8120 10900 8130 10940
rect 8170 10910 8320 10940
rect 8170 10900 8210 10910
rect 8120 10880 8210 10900
rect 7910 10810 8060 10840
rect 7910 10790 7950 10810
rect 7840 10770 7950 10790
rect 7350 10700 7380 10730
rect 7460 10700 7490 10730
rect 7920 10720 7950 10770
rect 8030 10720 8060 10810
rect 8180 10720 8210 10880
rect 8290 10720 8320 10910
rect 7350 10670 7490 10700
rect 7350 10420 7380 10670
rect 7250 10410 7380 10420
rect 7250 10350 7270 10410
rect 7330 10350 7380 10410
rect 7250 10340 7380 10350
rect 7350 10290 7380 10340
rect 7460 10290 7490 10670
rect 7350 9760 7380 9790
rect 7460 9760 7490 9790
rect 9930 10930 9960 10960
rect 10040 10930 10070 10960
rect 10470 10930 10500 10960
rect 10580 10930 10610 10960
rect 10730 10930 10760 10960
rect 10840 10930 10870 10960
rect 11070 10930 11100 10960
rect 11180 10930 11210 10960
rect 11460 10930 11490 10960
rect 11570 10930 11600 10960
rect 11720 10930 11750 10960
rect 11830 10930 11860 10960
rect 12060 10930 12090 10960
rect 12170 10930 12200 10960
rect 12460 10930 12490 10960
rect 12570 10930 12600 10960
rect 12720 10930 12750 10960
rect 12830 10930 12860 10960
rect 13060 10930 13090 10960
rect 13170 10930 13200 10960
rect 9930 10710 9960 10730
rect 10040 10710 10070 10730
rect 9090 10670 9120 10700
rect 9350 10670 9380 10700
rect 9600 10670 9630 10700
rect 9930 10690 10070 10710
rect 9840 10680 10070 10690
rect 8710 10430 8740 10580
rect 8860 10540 8890 10580
rect 8790 10520 8890 10540
rect 8790 10480 8810 10520
rect 8850 10480 8890 10520
rect 8790 10460 8890 10480
rect 9840 10640 9860 10680
rect 9900 10640 9960 10680
rect 9840 10630 9960 10640
rect 8640 10410 8740 10430
rect 8640 10370 8660 10410
rect 8700 10370 8740 10410
rect 8640 10350 8740 10370
rect 8710 10300 8740 10350
rect 8860 10300 8890 10460
rect 9090 10420 9120 10470
rect 9350 10420 9380 10470
rect 9600 10420 9630 10470
rect 9020 10400 9120 10420
rect 9020 10360 9040 10400
rect 9080 10360 9120 10400
rect 9020 10340 9120 10360
rect 9280 10400 9380 10420
rect 9280 10360 9300 10400
rect 9340 10360 9380 10400
rect 9280 10340 9380 10360
rect 9530 10400 9630 10420
rect 9530 10360 9550 10400
rect 9590 10360 9630 10400
rect 9530 10340 9630 10360
rect 9090 10300 9120 10340
rect 9350 10300 9380 10340
rect 9600 10300 9630 10340
rect 9930 10290 9960 10630
rect 10040 10390 10070 10680
rect 10470 10410 10500 10530
rect 10410 10390 10500 10410
rect 10410 10350 10420 10390
rect 10460 10380 10500 10390
rect 10580 10380 10610 10530
rect 10730 10510 10760 10530
rect 10670 10490 10760 10510
rect 10670 10450 10680 10490
rect 10720 10480 10760 10490
rect 10840 10480 10870 10530
rect 10720 10450 10870 10480
rect 10670 10430 10760 10450
rect 10460 10350 10610 10380
rect 10410 10330 10500 10350
rect 10040 10290 10070 10330
rect 10470 10290 10500 10330
rect 10580 10290 10610 10350
rect 10730 10290 10760 10430
rect 10840 10290 10870 10450
rect 11070 10390 11100 10730
rect 11180 10390 11210 10730
rect 11460 10410 11490 10530
rect 11400 10390 11490 10410
rect 10980 10380 11100 10390
rect 10980 10340 11000 10380
rect 11040 10340 11100 10380
rect 10980 10330 11100 10340
rect 11400 10350 11410 10390
rect 11450 10380 11490 10390
rect 11570 10380 11600 10530
rect 11720 10510 11750 10530
rect 11660 10490 11750 10510
rect 11660 10450 11670 10490
rect 11710 10480 11750 10490
rect 11830 10480 11860 10530
rect 11710 10450 11860 10480
rect 11660 10430 11750 10450
rect 11450 10350 11600 10380
rect 11400 10330 11490 10350
rect 11070 10290 11100 10330
rect 11180 10290 11210 10330
rect 11460 10290 11490 10330
rect 11570 10290 11600 10350
rect 11720 10290 11750 10430
rect 11830 10290 11860 10450
rect 12060 10390 12090 10730
rect 12170 10390 12200 10730
rect 12460 10410 12490 10530
rect 12400 10390 12490 10410
rect 11970 10380 12090 10390
rect 11970 10340 11990 10380
rect 12030 10340 12090 10380
rect 11970 10330 12090 10340
rect 12400 10350 12410 10390
rect 12450 10380 12490 10390
rect 12570 10380 12600 10530
rect 12720 10510 12750 10530
rect 12660 10490 12750 10510
rect 12660 10450 12670 10490
rect 12710 10480 12750 10490
rect 12830 10480 12860 10530
rect 12710 10450 12860 10480
rect 12660 10430 12750 10450
rect 12450 10350 12600 10380
rect 12400 10330 12490 10350
rect 12060 10290 12090 10330
rect 12170 10290 12200 10330
rect 12460 10290 12490 10330
rect 12570 10290 12600 10350
rect 12720 10290 12750 10430
rect 12830 10290 12860 10450
rect 13060 10390 13090 10730
rect 12970 10380 13090 10390
rect 12970 10340 12990 10380
rect 13030 10340 13090 10380
rect 12970 10330 13090 10340
rect 13060 10290 13090 10330
rect 13170 10290 13200 10730
rect 13400 10650 13430 10680
rect 13630 10650 13660 10680
rect 13740 10650 13770 10680
rect 13970 10650 14000 10680
rect 14080 10650 14110 10680
rect 14190 10650 14220 10680
rect 14300 10650 14330 10680
rect 14530 10650 14560 10680
rect 14640 10650 14670 10680
rect 14750 10650 14780 10680
rect 14860 10650 14890 10680
rect 14970 10650 15000 10680
rect 15080 10650 15110 10680
rect 15190 10650 15220 10680
rect 15300 10650 15330 10680
rect 15590 10650 15620 10680
rect 15700 10650 15730 10680
rect 15810 10650 15840 10680
rect 15920 10650 15950 10680
rect 16030 10650 16060 10680
rect 16140 10650 16170 10680
rect 16250 10650 16280 10680
rect 16360 10650 16390 10680
rect 16470 10650 16500 10680
rect 16580 10650 16610 10680
rect 16690 10650 16720 10680
rect 16800 10650 16830 10680
rect 16910 10650 16940 10680
rect 17020 10650 17050 10680
rect 17130 10650 17160 10680
rect 17240 10650 17270 10680
rect 17540 10650 17570 10680
rect 17650 10650 17680 10680
rect 17760 10650 17790 10680
rect 17870 10650 17900 10680
rect 17980 10650 18010 10680
rect 18090 10650 18120 10680
rect 18200 10650 18230 10680
rect 18310 10650 18340 10680
rect 18420 10650 18450 10680
rect 18530 10650 18560 10680
rect 18640 10650 18670 10680
rect 18750 10650 18780 10680
rect 18860 10650 18890 10680
rect 18970 10650 19000 10680
rect 19080 10650 19110 10680
rect 19190 10650 19220 10680
rect 19300 10650 19330 10680
rect 19410 10650 19440 10680
rect 19520 10650 19550 10680
rect 19630 10650 19660 10680
rect 19740 10650 19770 10680
rect 19850 10650 19880 10680
rect 19960 10650 19990 10680
rect 20070 10650 20100 10680
rect 20180 10650 20210 10680
rect 20290 10650 20320 10680
rect 20400 10650 20430 10680
rect 20510 10650 20540 10680
rect 20620 10650 20650 10680
rect 20730 10650 20760 10680
rect 20840 10650 20870 10680
rect 20950 10650 20980 10680
rect 13400 10410 13430 10450
rect 13630 10410 13660 10450
rect 13740 10410 13770 10450
rect 13970 10410 14000 10450
rect 14080 10410 14110 10450
rect 14190 10410 14220 10450
rect 14300 10410 14330 10450
rect 14530 10410 14560 10450
rect 14640 10410 14670 10450
rect 14750 10410 14780 10450
rect 14860 10410 14890 10450
rect 14970 10410 15000 10450
rect 15080 10410 15110 10450
rect 15190 10410 15220 10450
rect 15300 10410 15330 10450
rect 15590 10410 15620 10450
rect 15700 10410 15730 10450
rect 15810 10410 15840 10450
rect 15920 10410 15950 10450
rect 16030 10410 16060 10450
rect 16140 10410 16170 10450
rect 16250 10410 16280 10450
rect 16360 10410 16390 10450
rect 16470 10410 16500 10450
rect 16580 10410 16610 10450
rect 16690 10410 16720 10450
rect 16800 10410 16830 10450
rect 16910 10410 16940 10450
rect 17020 10410 17050 10450
rect 17130 10410 17160 10450
rect 17240 10410 17270 10450
rect 17540 10410 17570 10450
rect 17650 10410 17680 10450
rect 17760 10410 17790 10450
rect 17870 10410 17900 10450
rect 17980 10410 18010 10450
rect 18090 10410 18120 10450
rect 18200 10410 18230 10450
rect 18310 10410 18340 10450
rect 18420 10410 18450 10450
rect 18530 10410 18560 10450
rect 18640 10410 18670 10450
rect 18750 10410 18780 10450
rect 18860 10410 18890 10450
rect 18970 10410 19000 10450
rect 19080 10410 19110 10450
rect 19190 10410 19220 10450
rect 19300 10410 19330 10450
rect 19410 10410 19440 10450
rect 19520 10410 19550 10450
rect 19630 10410 19660 10450
rect 19740 10410 19770 10450
rect 19850 10410 19880 10450
rect 19960 10410 19990 10450
rect 20070 10410 20100 10450
rect 20180 10410 20210 10450
rect 20290 10410 20320 10450
rect 20400 10410 20430 10450
rect 20510 10410 20540 10450
rect 20620 10410 20650 10450
rect 20730 10410 20760 10450
rect 20840 10410 20870 10450
rect 20950 10410 20980 10450
rect 13340 10390 13430 10410
rect 13340 10350 13350 10390
rect 13390 10350 13430 10390
rect 13340 10330 13430 10350
rect 13570 10390 13770 10410
rect 13570 10350 13580 10390
rect 13620 10370 13770 10390
rect 13620 10350 13660 10370
rect 13570 10330 13660 10350
rect 13400 10290 13430 10330
rect 13630 10290 13660 10330
rect 13740 10290 13770 10370
rect 13910 10390 14330 10410
rect 13910 10350 13920 10390
rect 13960 10370 14330 10390
rect 13960 10350 14000 10370
rect 13910 10330 14000 10350
rect 13970 10290 14000 10330
rect 14080 10290 14110 10370
rect 14190 10290 14220 10370
rect 14300 10290 14330 10370
rect 14470 10390 15330 10410
rect 14470 10350 14480 10390
rect 14520 10370 15330 10390
rect 14520 10350 14560 10370
rect 14470 10330 14560 10350
rect 14530 10290 14560 10330
rect 14640 10290 14670 10370
rect 14750 10290 14780 10370
rect 14860 10290 14890 10370
rect 14970 10290 15000 10370
rect 15080 10290 15110 10370
rect 15190 10290 15220 10370
rect 15300 10290 15330 10370
rect 15530 10390 17270 10410
rect 15530 10350 15540 10390
rect 15580 10370 17270 10390
rect 15580 10350 15620 10370
rect 15530 10330 15620 10350
rect 15590 10290 15620 10330
rect 15700 10290 15730 10370
rect 15810 10290 15840 10370
rect 15920 10290 15950 10370
rect 16030 10290 16060 10370
rect 16140 10290 16170 10370
rect 16250 10290 16280 10370
rect 16360 10290 16390 10370
rect 16470 10290 16500 10370
rect 16580 10290 16610 10370
rect 16690 10290 16720 10370
rect 16800 10290 16830 10370
rect 16910 10290 16940 10370
rect 17020 10290 17050 10370
rect 17130 10290 17160 10370
rect 17240 10290 17270 10370
rect 17470 10390 20980 10410
rect 17470 10350 17490 10390
rect 17530 10370 20980 10390
rect 17530 10350 17570 10370
rect 17470 10330 17570 10350
rect 17540 10290 17570 10330
rect 17650 10290 17680 10370
rect 17760 10290 17790 10370
rect 17870 10290 17900 10370
rect 17980 10290 18010 10370
rect 18090 10290 18120 10370
rect 18200 10290 18230 10370
rect 18310 10290 18340 10370
rect 18420 10290 18450 10370
rect 18530 10290 18560 10370
rect 18640 10290 18670 10370
rect 18750 10290 18780 10370
rect 18860 10290 18890 10370
rect 18970 10290 19000 10370
rect 19080 10290 19110 10370
rect 19190 10290 19220 10370
rect 19300 10290 19330 10370
rect 19410 10290 19440 10370
rect 19520 10290 19550 10370
rect 19630 10290 19660 10370
rect 19740 10290 19770 10370
rect 19850 10290 19880 10370
rect 19960 10290 19990 10370
rect 20070 10290 20100 10370
rect 20180 10290 20210 10370
rect 20290 10290 20320 10370
rect 20400 10290 20430 10370
rect 20510 10290 20540 10370
rect 20620 10290 20650 10370
rect 20730 10290 20760 10370
rect 20840 10290 20870 10370
rect 20950 10290 20980 10370
rect 8710 9770 8740 9800
rect 8860 9770 8890 9800
rect 9090 9770 9120 9800
rect 9350 9770 9380 9800
rect 9600 9770 9630 9800
rect 9930 9760 9960 9790
rect 10040 9760 10070 9790
rect 10470 9760 10500 9790
rect 10580 9760 10610 9790
rect 10730 9760 10760 9790
rect 10840 9760 10870 9790
rect 11070 9760 11100 9790
rect 11180 9760 11210 9790
rect 11460 9760 11490 9790
rect 11570 9760 11600 9790
rect 11720 9760 11750 9790
rect 11830 9760 11860 9790
rect 12060 9760 12090 9790
rect 12170 9760 12200 9790
rect 12460 9760 12490 9790
rect 12570 9760 12600 9790
rect 12720 9760 12750 9790
rect 12830 9760 12860 9790
rect 13060 9760 13090 9790
rect 13170 9760 13200 9790
rect 13400 9760 13430 9790
rect 13630 9760 13660 9790
rect 13740 9760 13770 9790
rect 13970 9760 14000 9790
rect 14080 9760 14110 9790
rect 14190 9760 14220 9790
rect 14300 9760 14330 9790
rect 14530 9760 14560 9790
rect 14640 9760 14670 9790
rect 14750 9760 14780 9790
rect 14860 9760 14890 9790
rect 14970 9760 15000 9790
rect 15080 9760 15110 9790
rect 15190 9760 15220 9790
rect 15300 9760 15330 9790
rect 15590 9760 15620 9790
rect 15700 9760 15730 9790
rect 15810 9760 15840 9790
rect 15920 9760 15950 9790
rect 16030 9760 16060 9790
rect 16140 9760 16170 9790
rect 16250 9760 16280 9790
rect 16360 9760 16390 9790
rect 16470 9760 16500 9790
rect 16580 9760 16610 9790
rect 16690 9760 16720 9790
rect 16800 9760 16830 9790
rect 16910 9760 16940 9790
rect 17020 9760 17050 9790
rect 17130 9760 17160 9790
rect 17240 9760 17270 9790
rect 17540 9760 17570 9790
rect 17650 9760 17680 9790
rect 17760 9760 17790 9790
rect 17870 9760 17900 9790
rect 17980 9760 18010 9790
rect 18090 9760 18120 9790
rect 18200 9760 18230 9790
rect 18310 9760 18340 9790
rect 18420 9760 18450 9790
rect 18530 9760 18560 9790
rect 18640 9760 18670 9790
rect 18750 9760 18780 9790
rect 18860 9760 18890 9790
rect 18970 9760 19000 9790
rect 19080 9760 19110 9790
rect 19190 9760 19220 9790
rect 19300 9760 19330 9790
rect 19410 9760 19440 9790
rect 19520 9760 19550 9790
rect 19630 9760 19660 9790
rect 19740 9760 19770 9790
rect 19850 9760 19880 9790
rect 19960 9760 19990 9790
rect 20070 9760 20100 9790
rect 20180 9760 20210 9790
rect 20290 9760 20320 9790
rect 20400 9760 20430 9790
rect 20510 9760 20540 9790
rect 20620 9760 20650 9790
rect 20730 9760 20760 9790
rect 20840 9760 20870 9790
rect 20950 9760 20980 9790
rect 7920 9690 7950 9720
rect 8030 9690 8060 9720
rect 8180 9690 8210 9720
rect 8290 9690 8320 9720
rect 13160 8630 13300 8640
rect 13160 8580 13220 8630
rect 13270 8580 13300 8630
rect 13160 8570 13300 8580
rect 13160 8370 13190 8570
rect 9970 8340 13190 8370
rect 9970 8260 10000 8340
rect 10080 8260 10110 8340
rect 10190 8260 10220 8340
rect 10300 8260 10330 8340
rect 10410 8260 10440 8340
rect 10520 8260 10550 8340
rect 10630 8260 10660 8340
rect 10740 8260 10770 8340
rect 10850 8260 10880 8340
rect 10960 8260 10990 8340
rect 11070 8260 11100 8340
rect 11180 8260 11210 8340
rect 11290 8260 11320 8340
rect 11400 8260 11430 8340
rect 11510 8260 11540 8340
rect 11620 8260 11650 8340
rect 11730 8260 11760 8340
rect 11840 8260 11870 8340
rect 11950 8260 11980 8340
rect 12060 8260 12090 8340
rect 12170 8260 12200 8340
rect 12280 8260 12310 8340
rect 12390 8260 12420 8340
rect 12500 8260 12530 8340
rect 12610 8260 12640 8340
rect 12720 8260 12750 8340
rect 12830 8260 12860 8340
rect 12940 8260 12970 8340
rect 13050 8260 13080 8340
rect 13160 8260 13190 8340
rect 13740 8360 17130 8370
rect 13740 8340 17050 8360
rect 13740 8260 13770 8340
rect 13850 8260 13880 8340
rect 13960 8260 13990 8340
rect 14070 8260 14100 8340
rect 14180 8260 14210 8340
rect 14290 8260 14320 8340
rect 14400 8260 14430 8340
rect 14510 8260 14540 8340
rect 14620 8260 14650 8340
rect 14730 8260 14760 8340
rect 14840 8260 14870 8340
rect 14950 8260 14980 8340
rect 15060 8260 15090 8340
rect 15170 8260 15200 8340
rect 15280 8260 15310 8340
rect 15390 8260 15420 8340
rect 15500 8260 15530 8340
rect 15610 8260 15640 8340
rect 15720 8260 15750 8340
rect 15830 8260 15860 8340
rect 15940 8260 15970 8340
rect 16050 8260 16080 8340
rect 16160 8260 16190 8340
rect 16270 8260 16300 8340
rect 16380 8260 16410 8340
rect 16490 8260 16520 8340
rect 16600 8260 16630 8340
rect 16710 8260 16740 8340
rect 16820 8260 16850 8340
rect 16930 8310 17050 8340
rect 17100 8310 17130 8360
rect 16930 8300 17130 8310
rect 16930 8260 16960 8300
rect 9970 7030 10000 7060
rect 10080 7030 10110 7060
rect 10190 7030 10220 7060
rect 10300 7030 10330 7060
rect 10410 7030 10440 7060
rect 10520 7030 10550 7060
rect 10630 7030 10660 7060
rect 10740 7030 10770 7060
rect 10850 7030 10880 7060
rect 10960 7030 10990 7060
rect 11070 7030 11100 7060
rect 11180 7030 11210 7060
rect 11290 7030 11320 7060
rect 11400 7030 11430 7060
rect 11510 7030 11540 7060
rect 11620 7030 11650 7060
rect 11730 7030 11760 7060
rect 11840 7030 11870 7060
rect 11950 7030 11980 7060
rect 12060 7030 12090 7060
rect 12170 7030 12200 7060
rect 12280 7030 12310 7060
rect 12390 7030 12420 7060
rect 12500 7030 12530 7060
rect 12610 7030 12640 7060
rect 12720 7030 12750 7060
rect 12830 7030 12860 7060
rect 12940 7030 12970 7060
rect 13050 7030 13080 7060
rect 13160 7030 13190 7060
rect 13740 7030 13770 7060
rect 13850 7030 13880 7060
rect 13960 7030 13990 7060
rect 14070 7030 14100 7060
rect 14180 7030 14210 7060
rect 14290 7030 14320 7060
rect 14400 7030 14430 7060
rect 14510 7030 14540 7060
rect 14620 7030 14650 7060
rect 14730 7030 14760 7060
rect 14840 7030 14870 7060
rect 14950 7030 14980 7060
rect 15060 7030 15090 7060
rect 15170 7030 15200 7060
rect 15280 7030 15310 7060
rect 15390 7030 15420 7060
rect 15500 7030 15530 7060
rect 15610 7030 15640 7060
rect 15720 7030 15750 7060
rect 15830 7030 15860 7060
rect 15940 7030 15970 7060
rect 16050 7030 16080 7060
rect 16160 7030 16190 7060
rect 16270 7030 16300 7060
rect 16380 7030 16410 7060
rect 16490 7030 16520 7060
rect 16600 7030 16630 7060
rect 16710 7030 16740 7060
rect 16820 7030 16850 7060
rect 16930 7030 16960 7060
rect 13700 5860 13730 5890
rect 13810 5860 13840 5890
rect 13920 5860 13950 5890
rect 14030 5860 14060 5890
rect 14140 5860 14170 5890
rect 14250 5860 14280 5890
rect 14360 5860 14390 5890
rect 14470 5860 14500 5890
rect 14580 5860 14610 5890
rect 14690 5860 14720 5890
rect 14800 5860 14830 5890
rect 14910 5860 14940 5890
rect 15020 5860 15050 5890
rect 15130 5860 15160 5890
rect 15240 5860 15270 5890
rect 15350 5860 15380 5890
rect 15460 5860 15490 5890
rect 15570 5860 15600 5890
rect 15680 5860 15710 5890
rect 15790 5860 15820 5890
rect 15900 5860 15930 5890
rect 16010 5860 16040 5890
rect 16120 5860 16150 5890
rect 16230 5860 16260 5890
rect 16340 5860 16370 5890
rect 16450 5860 16480 5890
rect 16560 5860 16590 5890
rect 16670 5860 16700 5890
rect 16780 5860 16810 5890
rect 16890 5860 16920 5890
rect 9940 5620 9970 5650
rect 10050 5620 10080 5650
rect 10160 5620 10190 5650
rect 10270 5620 10300 5650
rect 10380 5620 10410 5650
rect 10490 5620 10520 5650
rect 10600 5620 10630 5650
rect 10710 5620 10740 5650
rect 10820 5620 10850 5650
rect 10930 5620 10960 5650
rect 11040 5620 11070 5650
rect 11150 5620 11180 5650
rect 11260 5620 11290 5650
rect 11370 5620 11400 5650
rect 11480 5620 11510 5650
rect 11590 5620 11620 5650
rect 11700 5620 11730 5650
rect 11810 5620 11840 5650
rect 11920 5620 11950 5650
rect 12030 5620 12060 5650
rect 12140 5620 12170 5650
rect 12250 5620 12280 5650
rect 12360 5620 12390 5650
rect 12470 5620 12500 5650
rect 12580 5620 12610 5650
rect 12690 5620 12720 5650
rect 12800 5620 12830 5650
rect 12910 5620 12940 5650
rect 13020 5620 13050 5650
rect 13130 5620 13160 5650
rect 13700 4580 13730 4660
rect 13810 4580 13840 4660
rect 13920 4580 13950 4660
rect 14030 4580 14060 4660
rect 14140 4580 14170 4660
rect 14250 4580 14280 4660
rect 14360 4580 14390 4660
rect 14470 4580 14500 4660
rect 14580 4580 14610 4660
rect 14690 4580 14720 4660
rect 14800 4580 14830 4660
rect 14910 4580 14940 4660
rect 15020 4580 15050 4660
rect 15130 4580 15160 4660
rect 15240 4580 15270 4660
rect 15350 4580 15380 4660
rect 15460 4580 15490 4660
rect 15570 4580 15600 4660
rect 15680 4580 15710 4660
rect 15790 4580 15820 4660
rect 15900 4580 15930 4660
rect 16010 4580 16040 4660
rect 16120 4580 16150 4660
rect 16230 4580 16260 4660
rect 16340 4580 16370 4660
rect 16450 4580 16480 4660
rect 16560 4580 16590 4660
rect 16670 4580 16700 4660
rect 16780 4580 16810 4660
rect 16890 4580 16920 4660
rect 13700 4550 16920 4580
rect 16890 4480 16920 4550
rect 16890 4470 17030 4480
rect 16890 4420 16950 4470
rect 17000 4420 17030 4470
rect 9940 4340 9970 4420
rect 10050 4340 10080 4420
rect 10160 4340 10190 4420
rect 10270 4340 10300 4420
rect 10380 4340 10410 4420
rect 10490 4340 10520 4420
rect 10600 4340 10630 4420
rect 10710 4340 10740 4420
rect 10820 4340 10850 4420
rect 10930 4340 10960 4420
rect 11040 4340 11070 4420
rect 11150 4340 11180 4420
rect 11260 4340 11290 4420
rect 11370 4340 11400 4420
rect 11480 4340 11510 4420
rect 11590 4340 11620 4420
rect 11700 4340 11730 4420
rect 11810 4340 11840 4420
rect 11920 4340 11950 4420
rect 12030 4340 12060 4420
rect 12140 4340 12170 4420
rect 12250 4340 12280 4420
rect 12360 4340 12390 4420
rect 12470 4340 12500 4420
rect 12580 4340 12610 4420
rect 12690 4340 12720 4420
rect 12800 4340 12830 4420
rect 12910 4340 12940 4420
rect 13020 4340 13050 4420
rect 13130 4340 13160 4420
rect 16890 4410 17030 4420
rect 9940 4310 13160 4340
rect 13130 4170 13160 4310
rect 13130 4150 13270 4170
rect 13130 4090 13180 4150
rect 13250 4090 13270 4150
rect 13700 4140 13730 4170
rect 13810 4140 13840 4170
rect 13920 4140 13950 4170
rect 14030 4140 14060 4170
rect 14140 4140 14170 4170
rect 14250 4140 14280 4170
rect 14360 4140 14390 4170
rect 14470 4140 14500 4170
rect 14580 4140 14610 4170
rect 14690 4140 14720 4170
rect 14800 4140 14830 4170
rect 14910 4140 14940 4170
rect 15020 4140 15050 4170
rect 15130 4140 15160 4170
rect 15240 4140 15270 4170
rect 15350 4140 15380 4170
rect 15460 4140 15490 4170
rect 15570 4140 15600 4170
rect 15680 4140 15710 4170
rect 15790 4140 15820 4170
rect 15900 4140 15930 4170
rect 16010 4140 16040 4170
rect 16120 4140 16150 4170
rect 16230 4140 16260 4170
rect 16340 4140 16370 4170
rect 16450 4140 16480 4170
rect 16560 4140 16590 4170
rect 16670 4140 16700 4170
rect 16780 4140 16810 4170
rect 16890 4140 16920 4170
rect 13130 4070 13270 4090
rect 13130 3960 13270 3980
rect 13130 3900 13180 3960
rect 13250 3900 13270 3960
rect 13130 3880 13270 3900
rect 9940 3810 9970 3840
rect 10050 3810 10080 3840
rect 10160 3810 10190 3840
rect 10270 3810 10300 3840
rect 10380 3810 10410 3840
rect 10490 3810 10520 3840
rect 10600 3810 10630 3840
rect 10710 3810 10740 3840
rect 10820 3810 10850 3840
rect 10930 3810 10960 3840
rect 11040 3810 11070 3840
rect 11150 3810 11180 3840
rect 11260 3810 11290 3840
rect 11370 3810 11400 3840
rect 11480 3810 11510 3840
rect 11590 3810 11620 3840
rect 11700 3810 11730 3840
rect 11810 3810 11840 3840
rect 11920 3810 11950 3840
rect 12030 3810 12060 3840
rect 12140 3810 12170 3840
rect 12250 3810 12280 3840
rect 12360 3810 12390 3840
rect 12470 3810 12500 3840
rect 12580 3810 12610 3840
rect 12690 3810 12720 3840
rect 12800 3810 12830 3840
rect 12910 3810 12940 3840
rect 13020 3810 13050 3840
rect 13130 3810 13160 3880
rect 13700 3510 13730 3540
rect 13810 3510 13840 3540
rect 13920 3510 13950 3540
rect 14030 3510 14060 3540
rect 14140 3510 14170 3540
rect 14250 3510 14280 3540
rect 14360 3510 14390 3540
rect 14470 3510 14500 3540
rect 14580 3510 14610 3540
rect 14690 3510 14720 3540
rect 14800 3510 14830 3540
rect 14910 3510 14940 3540
rect 15020 3510 15050 3540
rect 15130 3510 15160 3540
rect 15240 3510 15270 3540
rect 15350 3510 15380 3540
rect 15460 3510 15490 3540
rect 15570 3510 15600 3540
rect 15680 3510 15710 3540
rect 15790 3510 15820 3540
rect 15900 3510 15930 3540
rect 16010 3510 16040 3540
rect 16120 3510 16150 3540
rect 16230 3510 16260 3540
rect 16340 3510 16370 3540
rect 16450 3510 16480 3540
rect 16560 3510 16590 3540
rect 16670 3510 16700 3540
rect 16780 3510 16810 3540
rect 16890 3510 16920 3540
rect 13700 3480 16920 3510
rect 16890 3250 16920 3480
rect 16890 3240 17020 3250
rect 9940 3180 9970 3210
rect 10050 3180 10080 3210
rect 10160 3180 10190 3210
rect 10270 3180 10300 3210
rect 10380 3180 10410 3210
rect 10490 3180 10520 3210
rect 10600 3180 10630 3210
rect 10710 3180 10740 3210
rect 10820 3180 10850 3210
rect 10930 3180 10960 3210
rect 11040 3180 11070 3210
rect 11150 3180 11180 3210
rect 11260 3180 11290 3210
rect 11370 3180 11400 3210
rect 11480 3180 11510 3210
rect 11590 3180 11620 3210
rect 11700 3180 11730 3210
rect 11810 3180 11840 3210
rect 11920 3180 11950 3210
rect 12030 3180 12060 3210
rect 12140 3180 12170 3210
rect 12250 3180 12280 3210
rect 12360 3180 12390 3210
rect 12470 3180 12500 3210
rect 12580 3180 12610 3210
rect 12690 3180 12720 3210
rect 12800 3180 12830 3210
rect 12910 3180 12940 3210
rect 13020 3180 13050 3210
rect 13130 3180 13160 3210
rect 16890 3190 16950 3240
rect 17000 3190 17020 3240
rect 16890 3180 17020 3190
rect 9940 3150 13160 3180
rect 25700 2760 25790 2790
rect 25700 2720 25720 2760
rect 25770 2720 25790 2760
rect 25700 2700 25790 2720
rect 24320 2670 24350 2700
rect 25350 2670 25790 2700
rect 25700 2640 25790 2670
rect 25700 2600 25720 2640
rect 25770 2600 25790 2640
rect 25700 2590 25790 2600
rect 24320 2560 24350 2590
rect 25350 2560 25790 2590
rect 25700 2520 25790 2560
rect 25700 2480 25720 2520
rect 25770 2480 25790 2520
rect 24320 2450 24350 2480
rect 25350 2450 25790 2480
rect 25700 2400 25790 2450
rect 25700 2370 25720 2400
rect 24320 2340 24350 2370
rect 25350 2360 25720 2370
rect 25770 2360 25790 2400
rect 25350 2340 25790 2360
rect 25700 2280 25790 2340
rect 25700 2260 25720 2280
rect 24320 2230 24350 2260
rect 25350 2240 25720 2260
rect 25770 2240 25790 2280
rect 25350 2230 25790 2240
rect 25700 2160 25790 2230
rect 25700 2150 25720 2160
rect 24320 2120 24350 2150
rect 25350 2120 25720 2150
rect 25770 2120 25790 2160
rect 25700 2060 25790 2120
rect 13150 1680 13280 1690
rect 13150 1630 13210 1680
rect 13260 1630 13280 1680
rect 13150 1620 13280 1630
rect 13150 1390 13180 1620
rect 9960 1360 13180 1390
rect 9960 1330 9990 1360
rect 10070 1330 10100 1360
rect 10180 1330 10210 1360
rect 10290 1330 10320 1360
rect 10400 1330 10430 1360
rect 10510 1330 10540 1360
rect 10620 1330 10650 1360
rect 10730 1330 10760 1360
rect 10840 1330 10870 1360
rect 10950 1330 10980 1360
rect 11060 1330 11090 1360
rect 11170 1330 11200 1360
rect 11280 1330 11310 1360
rect 11390 1330 11420 1360
rect 11500 1330 11530 1360
rect 11610 1330 11640 1360
rect 11720 1330 11750 1360
rect 11830 1330 11860 1360
rect 11940 1330 11970 1360
rect 12050 1330 12080 1360
rect 12160 1330 12190 1360
rect 12270 1330 12300 1360
rect 12380 1330 12410 1360
rect 12490 1330 12520 1360
rect 12600 1330 12630 1360
rect 12710 1330 12740 1360
rect 12820 1330 12850 1360
rect 12930 1330 12960 1360
rect 13040 1330 13070 1360
rect 13150 1330 13180 1360
rect 13700 1420 17130 1430
rect 13700 1400 17060 1420
rect 13700 1320 13730 1400
rect 13810 1320 13840 1400
rect 13920 1320 13950 1400
rect 14030 1320 14060 1400
rect 14140 1320 14170 1400
rect 14250 1320 14280 1400
rect 14360 1320 14390 1400
rect 14470 1320 14500 1400
rect 14580 1320 14610 1400
rect 14690 1320 14720 1400
rect 14800 1320 14830 1400
rect 14910 1320 14940 1400
rect 15020 1320 15050 1400
rect 15130 1320 15160 1400
rect 15240 1320 15270 1400
rect 15350 1320 15380 1400
rect 15460 1320 15490 1400
rect 15570 1320 15600 1400
rect 15680 1320 15710 1400
rect 15790 1320 15820 1400
rect 15900 1320 15930 1400
rect 16010 1320 16040 1400
rect 16120 1320 16150 1400
rect 16230 1320 16260 1400
rect 16340 1320 16370 1400
rect 16450 1320 16480 1400
rect 16560 1320 16590 1400
rect 16670 1320 16700 1400
rect 16780 1320 16810 1400
rect 16890 1370 17060 1400
rect 17110 1370 17130 1420
rect 16890 1360 17130 1370
rect 16890 1320 16920 1360
rect 9960 700 9990 730
rect 10070 700 10100 730
rect 10180 700 10210 730
rect 10290 700 10320 730
rect 10400 700 10430 730
rect 10510 700 10540 730
rect 10620 700 10650 730
rect 10730 700 10760 730
rect 10840 700 10870 730
rect 10950 700 10980 730
rect 11060 700 11090 730
rect 11170 700 11200 730
rect 11280 700 11310 730
rect 11390 700 11420 730
rect 11500 700 11530 730
rect 11610 700 11640 730
rect 11720 700 11750 730
rect 11830 700 11860 730
rect 11940 700 11970 730
rect 12050 700 12080 730
rect 12160 700 12190 730
rect 12270 700 12300 730
rect 12380 700 12410 730
rect 12490 700 12520 730
rect 12600 700 12630 730
rect 12710 700 12740 730
rect 12820 700 12850 730
rect 12930 700 12960 730
rect 13040 700 13070 730
rect 13150 700 13180 730
rect 13700 690 13730 720
rect 13810 690 13840 720
rect 13920 690 13950 720
rect 14030 690 14060 720
rect 14140 690 14170 720
rect 14250 690 14280 720
rect 14360 690 14390 720
rect 14470 690 14500 720
rect 14580 690 14610 720
rect 14690 690 14720 720
rect 14800 690 14830 720
rect 14910 690 14940 720
rect 15020 690 15050 720
rect 15130 690 15160 720
rect 15240 690 15270 720
rect 15350 690 15380 720
rect 15460 690 15490 720
rect 15570 690 15600 720
rect 15680 690 15710 720
rect 15790 690 15820 720
rect 15900 690 15930 720
rect 16010 690 16040 720
rect 16120 690 16150 720
rect 16230 690 16260 720
rect 16340 690 16370 720
rect 16450 690 16480 720
rect 16560 690 16590 720
rect 16670 690 16700 720
rect 16780 690 16810 720
rect 16890 690 16920 720
<< polycont >>
rect 23470 42280 23510 42320
rect 2789 42010 2829 42050
rect 22070 42070 22130 42130
rect 22590 42060 22630 42100
rect 23500 42170 23540 42210
rect 23110 42100 23150 42140
rect 23000 41990 23040 42030
rect 21850 41930 21890 41970
rect 2679 41580 2719 41620
rect 2899 41540 2939 41580
rect 23000 41870 23040 41910
rect 22590 41760 22630 41800
rect 23110 41760 23150 41800
rect 23500 41720 23540 41760
rect 5969 41240 6009 41280
rect 6199 41240 6239 41280
rect 6539 41240 6579 41280
rect 7099 41240 7139 41280
rect 8159 41240 8199 41280
rect 2989 40900 3029 40940
rect 3469 40950 3509 40990
rect 5359 40940 5399 40980
rect 2999 40620 3039 40660
rect 6369 39920 6409 39960
rect 2759 39650 2799 39690
rect 3339 39660 3379 39700
rect 5359 39660 5399 39700
rect 3760 34940 3810 34990
rect 4560 34930 4620 35000
rect 5420 34820 5470 34870
rect 6340 34810 6380 34850
rect 6720 34810 6760 34850
rect 7300 34800 7340 34840
rect 7680 34800 7720 34840
rect 8060 34800 8100 34840
rect 8440 34800 8480 34840
rect 9060 34910 9100 34950
rect 8800 34800 8840 34840
rect 9380 34800 9420 34840
rect 9760 34800 9800 34840
rect 10140 34800 10180 34840
rect 10520 34800 10560 34840
rect 15460 36070 15500 36110
rect 15570 35570 15640 35630
rect 16450 35430 16510 35490
rect 17580 35450 17620 35490
rect 17720 35450 17760 35490
rect 18040 35450 18080 35490
rect 18520 35450 18560 35490
rect 18660 35450 18700 35490
rect 18980 35450 19020 35490
rect 17870 35160 17910 35200
rect 19770 35450 19810 35490
rect 20020 35480 20060 35520
rect 17470 34860 17510 34900
rect 18410 34860 18450 34900
rect 18700 34860 18740 34900
rect 21430 35450 21470 35490
rect 22540 35450 22580 35490
rect 22680 35450 22720 35490
rect 23000 35450 23040 35490
rect 23480 35450 23520 35490
rect 23620 35450 23660 35490
rect 23940 35450 23980 35490
rect 19320 34910 19360 34950
rect 20920 34900 20980 34960
rect 19750 34750 19810 34810
rect 20020 34770 20060 34810
rect 19770 34620 19810 34660
rect 17690 34320 17730 34360
rect 18040 34320 18080 34360
rect 22830 35160 22870 35200
rect 24730 35450 24770 35490
rect 24980 35480 25020 35520
rect 22430 34860 22470 34900
rect 23370 34860 23410 34900
rect 23660 34860 23700 34900
rect 24280 34910 24320 34950
rect 24710 34750 24770 34810
rect 24980 34770 25020 34810
rect 24730 34620 24770 34660
rect 18630 34320 18670 34360
rect 18980 34320 19020 34360
rect 22650 34320 22690 34360
rect 23000 34320 23040 34360
rect 23590 34320 23630 34360
rect 23940 34320 23980 34360
rect 7180 34150 7220 34190
rect 14118 32340 14158 32380
rect 14008 31900 14048 31940
rect 14228 31850 14268 31890
rect 16450 31390 16510 31450
rect 17580 31390 17620 31430
rect 17720 31390 17760 31430
rect 18040 31390 18080 31430
rect 18520 31390 18560 31430
rect 18660 31390 18700 31430
rect 18980 31390 19020 31430
rect 14118 31270 14158 31310
rect 2160 30690 2210 30740
rect 2960 30680 3020 30740
rect 3820 30560 3860 30600
rect 4680 30560 4730 30610
rect 6400 30660 6440 30700
rect 6780 30660 6820 30700
rect 5540 30560 5590 30610
rect 7360 30650 7400 30690
rect 7740 30650 7780 30690
rect 8120 30650 8160 30690
rect 8500 30650 8540 30690
rect 9120 30760 9160 30800
rect 8860 30650 8900 30690
rect 9440 30650 9480 30690
rect 9820 30650 9860 30690
rect 10200 30650 10240 30690
rect 10580 30650 10620 30690
rect 10960 30650 11000 30690
rect 17870 31100 17910 31140
rect 20030 31390 20070 31430
rect 20280 31400 20320 31440
rect 17470 30800 17510 30840
rect 18410 30800 18450 30840
rect 18700 30800 18740 30840
rect 19320 30850 19360 30890
rect 21490 31380 21530 31420
rect 22600 31380 22640 31420
rect 22740 31380 22780 31420
rect 23060 31380 23100 31420
rect 23540 31380 23580 31420
rect 23680 31380 23720 31420
rect 24000 31380 24040 31420
rect 19580 30850 19620 30890
rect 20980 30840 21040 30900
rect 20010 30690 20070 30750
rect 20280 30710 20320 30750
rect 20030 30560 20070 30600
rect 17690 30260 17730 30300
rect 18040 30260 18080 30300
rect 22890 31090 22930 31130
rect 24990 31380 25030 31420
rect 25240 31410 25280 31450
rect 22490 30790 22530 30830
rect 23430 30790 23470 30830
rect 23720 30790 23760 30830
rect 24340 30840 24380 30880
rect 24600 30840 24640 30880
rect 24970 30680 25030 30740
rect 25240 30700 25280 30740
rect 24990 30550 25030 30590
rect 18630 30260 18670 30300
rect 18980 30260 19020 30300
rect 22710 30250 22750 30290
rect 23060 30250 23100 30290
rect 23650 30250 23690 30290
rect 24000 30250 24040 30290
rect 7240 30000 7280 30040
rect 7290 25130 7350 25190
rect 7820 25500 7880 25560
rect 8500 24900 8540 24940
rect 8880 24900 8920 24940
rect 9220 24910 9260 24950
rect 8650 24820 8690 24860
rect 9680 25910 9720 25950
rect 9940 25910 9980 25950
rect 9680 25020 9720 25060
rect 9580 24900 9620 24940
rect 9940 25020 9980 25060
rect 9840 24800 9880 24840
rect 10160 24910 10200 24950
rect 10670 25910 10710 25950
rect 10930 25910 10970 25950
rect 10670 25020 10710 25060
rect 10570 24900 10610 24940
rect 10930 25020 10970 25060
rect 11150 24910 11190 24950
rect 10830 24800 10870 24840
rect 11670 25910 11710 25950
rect 11930 25910 11970 25950
rect 11670 25020 11710 25060
rect 11570 24900 11610 24940
rect 11930 25020 11970 25060
rect 11830 24800 11870 24840
rect 12150 24910 12190 24950
rect 12530 24910 12570 24950
rect 13230 25890 13270 25930
rect 13570 25890 13610 25930
rect 13790 25890 13830 25930
rect 14130 25910 14170 25950
rect 14350 25910 14390 25950
rect 14570 25910 14610 25950
rect 14790 25910 14830 25950
rect 15190 25910 15230 25950
rect 15410 25910 15450 25950
rect 15630 25910 15670 25950
rect 15850 25910 15890 25950
rect 16070 25910 16110 25950
rect 16290 25910 16330 25950
rect 16510 25910 16550 25950
rect 16730 25910 16770 25950
rect 17140 25910 17180 25950
rect 17360 25910 17400 25950
rect 17580 25910 17620 25950
rect 17800 25910 17840 25950
rect 18020 25910 18060 25950
rect 18240 25910 18280 25950
rect 18460 25910 18500 25950
rect 18680 25910 18720 25950
rect 18900 25910 18940 25950
rect 19120 25910 19160 25950
rect 19340 25910 19380 25950
rect 19560 25910 19600 25950
rect 19780 25910 19820 25950
rect 20000 25910 20040 25950
rect 20220 25910 20260 25950
rect 20440 25910 20480 25950
rect 13230 25000 13270 25040
rect 12900 24900 12940 24940
rect 13130 24900 13170 24940
rect 13570 25000 13610 25040
rect 13470 24900 13510 24940
rect 13790 25000 13830 25040
rect 14130 25020 14170 25060
rect 14030 24900 14070 24940
rect 14350 25020 14390 25060
rect 14570 25020 14610 25060
rect 14790 25020 14830 25060
rect 15190 25020 15230 25060
rect 15090 24900 15130 24940
rect 15410 25020 15450 25060
rect 15630 25020 15670 25060
rect 15850 25020 15890 25060
rect 16070 25020 16110 25060
rect 16290 25020 16330 25060
rect 16510 25020 16550 25060
rect 16730 25020 16770 25060
rect 17140 25020 17180 25060
rect 17040 24900 17080 24940
rect 17360 25020 17400 25060
rect 17580 25020 17620 25060
rect 17800 25020 17840 25060
rect 18020 25020 18060 25060
rect 18240 25020 18280 25060
rect 18460 25020 18500 25060
rect 18680 25020 18720 25060
rect 18900 25020 18940 25060
rect 19120 25020 19160 25060
rect 19340 25020 19380 25060
rect 19560 25020 19600 25060
rect 19780 25020 19820 25060
rect 20000 25020 20040 25060
rect 20220 25020 20260 25060
rect 20440 25020 20480 25060
rect 7380 22640 7420 22680
rect 7640 22730 7680 22770
rect 7480 22520 7520 22560
rect 7960 22630 8000 22670
rect 7740 22520 7780 22560
rect 7480 21660 7520 21700
rect 7740 21640 7780 21680
rect 8650 22710 8690 22750
rect 8500 22630 8540 22670
rect 8880 22630 8920 22670
rect 9220 22640 9280 22700
rect 9580 22630 9620 22670
rect 9840 22730 9880 22770
rect 9680 22510 9720 22550
rect 10160 22620 10200 22660
rect 9940 22510 9980 22550
rect 9680 21630 9720 21670
rect 9940 21630 9980 21670
rect 10570 22630 10610 22670
rect 10830 22730 10870 22770
rect 10670 22510 10710 22550
rect 11150 22620 11190 22660
rect 10930 22510 10970 22550
rect 10670 21630 10710 21670
rect 10930 21630 10970 21670
rect 11570 22630 11610 22670
rect 11830 22730 11870 22770
rect 11670 22510 11710 22550
rect 12150 22620 12190 22660
rect 11930 22510 11970 22550
rect 11670 21630 11710 21670
rect 11930 21630 11970 21670
rect 12530 22620 12570 22660
rect 12900 22630 12940 22670
rect 13130 22630 13170 22670
rect 13470 22630 13510 22670
rect 13230 22530 13270 22570
rect 13570 22530 13610 22570
rect 14030 22630 14070 22670
rect 13790 22530 13830 22570
rect 14130 22510 14170 22550
rect 14350 22510 14390 22550
rect 14570 22510 14610 22550
rect 15090 22630 15130 22670
rect 14790 22510 14830 22550
rect 15190 22510 15230 22550
rect 15410 22510 15450 22550
rect 15630 22510 15670 22550
rect 15850 22510 15890 22550
rect 16070 22510 16110 22550
rect 16290 22510 16330 22550
rect 16510 22510 16550 22550
rect 17040 22630 17080 22670
rect 16730 22510 16770 22550
rect 17140 22510 17180 22550
rect 17360 22510 17400 22550
rect 17580 22510 17620 22550
rect 17800 22510 17840 22550
rect 18020 22510 18060 22550
rect 18240 22510 18280 22550
rect 18460 22510 18500 22550
rect 18680 22510 18720 22550
rect 18900 22510 18940 22550
rect 19120 22510 19160 22550
rect 19340 22510 19380 22550
rect 19560 22510 19600 22550
rect 19780 22510 19820 22550
rect 20000 22510 20040 22550
rect 20220 22510 20260 22550
rect 20440 22510 20480 22550
rect 13230 21640 13270 21680
rect 13570 21640 13610 21680
rect 13790 21640 13830 21680
rect 14130 21620 14170 21660
rect 14350 21620 14390 21660
rect 14570 21620 14610 21660
rect 14790 21620 14830 21660
rect 15190 21620 15230 21660
rect 15410 21620 15450 21660
rect 15630 21620 15670 21660
rect 15850 21620 15890 21660
rect 16070 21620 16110 21660
rect 16290 21620 16330 21660
rect 16510 21620 16550 21660
rect 16730 21620 16770 21660
rect 17140 21620 17180 21660
rect 17360 21620 17400 21660
rect 17580 21620 17620 21660
rect 17800 21620 17840 21660
rect 18020 21620 18060 21660
rect 18240 21620 18280 21660
rect 18460 21620 18500 21660
rect 18680 21620 18720 21660
rect 18900 21620 18940 21660
rect 19120 21620 19160 21660
rect 19340 21620 19380 21660
rect 19560 21620 19600 21660
rect 19780 21620 19820 21660
rect 20000 21620 20040 21660
rect 20220 21620 20260 21660
rect 20440 21620 20480 21660
rect 7400 19270 7440 19310
rect 7400 18390 7440 18430
rect 7300 18130 7340 18170
rect 7560 18240 7600 18280
rect 7970 18240 8010 18280
rect 8500 18310 8540 18350
rect 8880 18310 8920 18350
rect 8650 18230 8690 18270
rect 9220 18270 9280 18330
rect 9680 19320 9720 19360
rect 9940 19320 9980 19360
rect 9680 18430 9720 18470
rect 9580 18310 9620 18350
rect 9940 18430 9980 18470
rect 9840 18210 9880 18250
rect 10160 18320 10200 18360
rect 10670 19320 10710 19360
rect 10930 19320 10970 19360
rect 10670 18430 10710 18470
rect 10570 18310 10610 18350
rect 10930 18430 10970 18470
rect 10830 18210 10870 18250
rect 11150 18320 11190 18360
rect 11670 19310 11710 19350
rect 11930 19310 11970 19350
rect 11670 18420 11710 18460
rect 11570 18310 11610 18350
rect 11930 18420 11970 18460
rect 11830 18210 11870 18250
rect 12150 18320 12190 18360
rect 12530 18320 12570 18360
rect 13230 19300 13270 19340
rect 13570 19300 13610 19340
rect 13790 19300 13830 19340
rect 14130 19320 14170 19360
rect 14350 19320 14390 19360
rect 14570 19320 14610 19360
rect 14790 19320 14830 19360
rect 15190 19320 15230 19360
rect 15410 19320 15450 19360
rect 15630 19320 15670 19360
rect 15850 19320 15890 19360
rect 16070 19320 16110 19360
rect 16290 19320 16330 19360
rect 16510 19320 16550 19360
rect 16730 19320 16770 19360
rect 17140 19320 17180 19360
rect 17360 19320 17400 19360
rect 17580 19320 17620 19360
rect 17800 19320 17840 19360
rect 18020 19320 18060 19360
rect 18240 19320 18280 19360
rect 18460 19320 18500 19360
rect 18680 19320 18720 19360
rect 18900 19320 18940 19360
rect 19120 19320 19160 19360
rect 19340 19320 19380 19360
rect 19560 19320 19600 19360
rect 19780 19320 19820 19360
rect 20000 19320 20040 19360
rect 20220 19320 20260 19360
rect 20440 19320 20480 19360
rect 13230 18410 13270 18450
rect 12900 18310 12940 18350
rect 13130 18310 13170 18350
rect 13570 18410 13610 18450
rect 13470 18310 13510 18350
rect 13790 18410 13830 18450
rect 14130 18430 14170 18470
rect 14030 18310 14070 18350
rect 14350 18430 14390 18470
rect 14570 18430 14610 18470
rect 14790 18430 14830 18470
rect 15190 18430 15230 18470
rect 15090 18310 15130 18350
rect 15410 18430 15450 18470
rect 15630 18430 15670 18470
rect 15850 18430 15890 18470
rect 16070 18430 16110 18470
rect 16290 18430 16330 18470
rect 16510 18430 16550 18470
rect 16730 18430 16770 18470
rect 17140 18430 17180 18470
rect 17040 18310 17080 18350
rect 17360 18430 17400 18470
rect 17580 18430 17620 18470
rect 17800 18430 17840 18470
rect 18020 18430 18060 18470
rect 18240 18430 18280 18470
rect 18460 18430 18500 18470
rect 18680 18430 18720 18470
rect 18900 18430 18940 18470
rect 19120 18430 19160 18470
rect 19340 18430 19380 18470
rect 19560 18430 19600 18470
rect 19780 18430 19820 18470
rect 20000 18430 20040 18470
rect 20220 18430 20260 18470
rect 20440 18430 20480 18470
rect 9750 15050 9810 15110
rect 10280 14960 10350 15020
rect 10580 15070 10620 15110
rect 10900 14960 10940 15000
rect 11310 14970 11350 15010
rect 11570 15070 11610 15110
rect 11890 14960 11930 15000
rect 12310 14970 12350 15010
rect 12570 15070 12610 15110
rect 12890 14960 12930 15000
rect 13260 14970 13300 15010
rect 13490 14970 13530 15010
rect 13830 14970 13870 15010
rect 14390 14970 14430 15010
rect 15450 14970 15490 15010
rect 17400 14970 17440 15010
rect 7270 12650 7330 12710
rect 7820 12660 7860 12700
rect 8570 12650 8610 12690
rect 8080 12560 8120 12600
rect 8950 12660 8990 12700
rect 9210 12660 9250 12700
rect 9460 12660 9500 12700
rect 9860 12670 9900 12710
rect 10420 12660 10460 12700
rect 8720 12540 8760 12580
rect 11000 12670 11040 12710
rect 11410 12660 11450 12700
rect 10680 12560 10720 12600
rect 11990 12670 12030 12710
rect 12410 12660 12450 12700
rect 11670 12560 11710 12600
rect 12990 12670 13030 12710
rect 13360 12660 13400 12700
rect 12670 12560 12710 12600
rect 13590 12660 13630 12700
rect 13930 12660 13970 12700
rect 14490 12660 14530 12700
rect 15550 12660 15590 12700
rect 17500 12660 17540 12700
rect 7850 10790 7910 10850
rect 8130 10900 8170 10940
rect 7270 10350 7330 10410
rect 8810 10480 8850 10520
rect 9860 10640 9900 10680
rect 8660 10370 8700 10410
rect 9040 10360 9080 10400
rect 9300 10360 9340 10400
rect 9550 10360 9590 10400
rect 10420 10350 10460 10390
rect 10680 10450 10720 10490
rect 11000 10340 11040 10380
rect 11410 10350 11450 10390
rect 11670 10450 11710 10490
rect 11990 10340 12030 10380
rect 12410 10350 12450 10390
rect 12670 10450 12710 10490
rect 12990 10340 13030 10380
rect 13350 10350 13390 10390
rect 13580 10350 13620 10390
rect 13920 10350 13960 10390
rect 14480 10350 14520 10390
rect 15540 10350 15580 10390
rect 17490 10350 17530 10390
rect 13220 8580 13270 8630
rect 17050 8310 17100 8360
rect 16950 4420 17000 4470
rect 13180 4090 13250 4150
rect 13180 3900 13250 3960
rect 16950 3190 17000 3240
rect 25720 2720 25770 2760
rect 25720 2600 25770 2640
rect 25720 2480 25770 2520
rect 25720 2360 25770 2400
rect 25720 2240 25770 2280
rect 25720 2120 25770 2160
rect 13210 1630 13260 1680
rect 17060 1370 17110 1420
<< locali >>
rect 21790 43350 23630 43360
rect 21790 43280 21830 43350
rect 21890 43280 21930 43350
rect 21990 43280 22030 43350
rect 22090 43280 22130 43350
rect 22190 43280 22230 43350
rect 22290 43280 22330 43350
rect 22390 43280 22430 43350
rect 22490 43280 22530 43350
rect 22590 43280 22630 43350
rect 22690 43280 22730 43350
rect 22790 43280 22830 43350
rect 22890 43280 22930 43350
rect 22990 43280 23030 43350
rect 23090 43280 23130 43350
rect 23190 43280 23230 43350
rect 23290 43280 23330 43350
rect 23390 43280 23430 43350
rect 23490 43280 23530 43350
rect 23590 43280 23630 43350
rect 21790 43270 23630 43280
rect 21720 42860 21780 42880
rect 21720 42200 21730 42860
rect 21770 42200 21780 42860
rect 2439 42160 2999 42170
rect 2439 42110 2469 42160
rect 2519 42110 2559 42160
rect 2609 42110 2649 42160
rect 2699 42110 2739 42160
rect 2789 42110 2829 42160
rect 2879 42110 2919 42160
rect 2969 42110 2999 42160
rect 2439 42100 2999 42110
rect 2439 41380 2499 42100
rect 2559 41900 2619 42100
rect 2769 42050 2849 42060
rect 2769 42010 2789 42050
rect 2829 42010 2849 42050
rect 2769 42000 2849 42010
rect 21720 42000 21780 42200
rect 21830 42860 21890 43270
rect 21830 42200 21840 42860
rect 21880 42200 21890 42860
rect 21830 42180 21890 42200
rect 21950 42860 22010 42880
rect 21950 42200 21960 42860
rect 22000 42200 22010 42860
rect 2559 41740 2569 41900
rect 2609 41740 2619 41900
rect 2559 41720 2619 41740
rect 2669 41900 2729 41920
rect 2669 41740 2679 41900
rect 2719 41740 2729 41900
rect 2669 41630 2729 41740
rect 2779 41900 2839 42000
rect 21610 41980 21780 42000
rect 5949 41970 9979 41980
rect 3390 41950 4329 41960
rect 2779 41740 2789 41900
rect 2829 41740 2839 41900
rect 2659 41620 2739 41630
rect 2659 41580 2679 41620
rect 2719 41580 2739 41620
rect 2659 41570 2739 41580
rect 2779 41510 2839 41740
rect 2889 41900 2949 41920
rect 2889 41740 2899 41900
rect 2939 41740 2949 41900
rect 3390 41900 3429 41950
rect 3479 41900 3519 41950
rect 3569 41900 3609 41950
rect 3659 41900 3699 41950
rect 3749 41900 3789 41950
rect 3839 41900 3879 41950
rect 3929 41900 3969 41950
rect 4019 41900 4059 41950
rect 4109 41900 4149 41950
rect 4199 41900 4239 41950
rect 4289 41900 4329 41950
rect 3390 41890 4329 41900
rect 4399 41950 5479 41960
rect 4399 41890 4579 41950
rect 4639 41890 5479 41950
rect 2889 41690 2949 41740
rect 3389 41800 3449 41890
rect 4399 41880 5479 41890
rect 5949 41910 6009 41970
rect 6069 41910 6119 41970
rect 6179 41910 6229 41970
rect 6289 41910 6339 41970
rect 6399 41910 6449 41970
rect 6509 41910 6559 41970
rect 6619 41910 6669 41970
rect 6729 41910 6779 41970
rect 6839 41910 6889 41970
rect 6949 41910 6999 41970
rect 7059 41910 7109 41970
rect 7169 41910 7219 41970
rect 7279 41910 7329 41970
rect 7389 41910 7439 41970
rect 7499 41910 7549 41970
rect 7609 41910 7659 41970
rect 7719 41910 7769 41970
rect 7829 41910 7879 41970
rect 7939 41910 7989 41970
rect 8049 41910 8099 41970
rect 8159 41910 8209 41970
rect 8269 41910 8319 41970
rect 8379 41910 8429 41970
rect 8489 41910 8539 41970
rect 8599 41910 8649 41970
rect 8709 41910 8759 41970
rect 8819 41910 8869 41970
rect 8929 41910 8979 41970
rect 9039 41910 9089 41970
rect 9149 41910 9199 41970
rect 9259 41910 9309 41970
rect 9369 41910 9419 41970
rect 9479 41910 9529 41970
rect 9589 41910 9639 41970
rect 9699 41910 9749 41970
rect 9809 41910 9859 41970
rect 9919 41910 9979 41970
rect 5949 41900 9979 41910
rect 21610 41920 21630 41980
rect 21700 41920 21780 41980
rect 21820 41970 21910 41980
rect 21950 41970 22010 42200
rect 22060 42860 22120 43270
rect 22320 43150 22420 43170
rect 22320 43090 22340 43150
rect 22400 43090 22640 43150
rect 22320 43070 22420 43090
rect 22060 42200 22070 42860
rect 22110 42200 22120 42860
rect 22060 42180 22120 42200
rect 22580 42870 22640 43090
rect 22580 42210 22590 42870
rect 22630 42210 22640 42870
rect 22580 42190 22640 42210
rect 22690 43040 23050 43090
rect 22690 42870 22750 43040
rect 22690 42210 22700 42870
rect 22740 42210 22750 42870
rect 22690 42190 22750 42210
rect 22880 42870 22940 42890
rect 22880 42210 22890 42870
rect 22930 42210 22940 42870
rect 22050 42130 22150 42140
rect 22050 42070 22070 42130
rect 22130 42070 22150 42130
rect 22050 42060 22150 42070
rect 22570 42100 22650 42110
rect 22570 42060 22590 42100
rect 22630 42060 22650 42100
rect 22570 42050 22650 42060
rect 22220 41970 22260 42030
rect 22580 41990 22630 42050
rect 22880 41990 22940 42210
rect 22990 42870 23050 43040
rect 22990 42210 23000 42870
rect 23040 42210 23050 42870
rect 22990 42190 23050 42210
rect 23100 42870 23160 43270
rect 23100 42210 23110 42870
rect 23150 42210 23160 42870
rect 23460 43160 23520 43180
rect 23460 42500 23470 43160
rect 23510 42500 23520 43160
rect 23460 42420 23520 42500
rect 23570 43160 23630 43270
rect 23570 42500 23580 43160
rect 23620 42500 23630 43160
rect 23570 42480 23630 42500
rect 23100 42190 23160 42210
rect 23280 42380 23520 42420
rect 23090 42140 23170 42150
rect 23090 42100 23110 42140
rect 23150 42100 23170 42140
rect 23090 42090 23170 42100
rect 22580 41970 22940 41990
rect 22980 42030 23060 42040
rect 23110 42030 23150 42090
rect 22980 41990 23000 42030
rect 23040 41990 23150 42030
rect 23280 41990 23330 42380
rect 23450 42320 23530 42330
rect 23450 42280 23470 42320
rect 23510 42280 23530 42320
rect 23450 42270 23530 42280
rect 23480 42210 23560 42220
rect 23480 42170 23500 42210
rect 23540 42170 23560 42210
rect 23480 42160 23560 42170
rect 22980 41980 23060 41990
rect 21820 41930 21850 41970
rect 21890 41930 22590 41970
rect 22630 41930 22940 41970
rect 21820 41920 21910 41930
rect 21610 41900 21780 41920
rect 3049 41690 3209 41700
rect 2889 41680 3209 41690
rect 2889 41640 3089 41680
rect 3169 41640 3209 41680
rect 2889 41630 3209 41640
rect 3049 41620 3209 41630
rect 2879 41580 2959 41590
rect 2879 41540 2899 41580
rect 2939 41540 2959 41580
rect 2879 41530 2959 41540
rect 2779 41470 2789 41510
rect 2829 41470 2839 41510
rect 2779 41450 2839 41470
rect 2439 41020 2449 41380
rect 2489 41020 2499 41380
rect 2439 41000 2499 41020
rect 2549 41380 2609 41400
rect 2549 41020 2559 41380
rect 2599 41020 2609 41380
rect 2549 40820 2609 41020
rect 2659 41380 2719 41400
rect 2659 41020 2669 41380
rect 2709 41020 2719 41380
rect 2659 41000 2719 41020
rect 2769 41380 2829 41400
rect 2769 41020 2779 41380
rect 2819 41020 2829 41380
rect 2769 41000 2829 41020
rect 2879 41380 2939 41400
rect 2879 41020 2889 41380
rect 2929 41020 2939 41380
rect 2879 41000 2939 41020
rect 2989 41380 3049 41400
rect 2989 41020 2999 41380
rect 3039 41020 3049 41380
rect 3389 41090 3399 41800
rect 3439 41090 3449 41800
rect 3389 41070 3449 41090
rect 3499 41800 3559 41820
rect 3499 41090 3509 41800
rect 3549 41090 3559 41800
rect 3499 41070 3559 41090
rect 3609 41800 3669 41820
rect 3609 41090 3619 41800
rect 3659 41090 3669 41800
rect 3609 41070 3669 41090
rect 3719 41800 3779 41820
rect 3719 41090 3729 41800
rect 3769 41090 3779 41800
rect 3719 41070 3779 41090
rect 3829 41800 3889 41820
rect 3829 41090 3839 41800
rect 3879 41090 3889 41800
rect 3829 41070 3889 41090
rect 3939 41800 3999 41820
rect 3939 41090 3949 41800
rect 3989 41090 3999 41800
rect 3939 41070 3999 41090
rect 4049 41800 4109 41820
rect 4049 41090 4059 41800
rect 4099 41090 4109 41800
rect 4049 41070 4109 41090
rect 4159 41800 4219 41820
rect 4159 41090 4169 41800
rect 4209 41090 4219 41800
rect 2989 41000 3049 41020
rect 3459 40990 3519 41010
rect 2979 40940 3039 40960
rect 2979 40900 2989 40940
rect 3029 40900 3039 40940
rect 3459 40950 3469 40990
rect 3509 40950 3519 40990
rect 3459 40930 3519 40950
rect 4159 40980 4219 41090
rect 4269 41800 4329 41820
rect 4269 41090 4279 41800
rect 4319 41090 4329 41800
rect 4269 41070 4329 41090
rect 4399 40980 4459 41880
rect 4159 40940 4459 40980
rect 4539 41790 4599 41880
rect 5949 41820 6009 41900
rect 4539 41080 4549 41790
rect 4589 41080 4599 41790
rect 2979 40870 3039 40900
rect 4539 40870 4599 41080
rect 2979 40830 4599 40870
rect 4649 41790 4709 41810
rect 4649 41080 4659 41790
rect 4699 41080 4709 41790
rect 2549 40770 2819 40820
rect 2759 40660 2819 40770
rect 2759 40620 2769 40660
rect 2809 40620 2819 40660
rect 2649 40540 2709 40560
rect 2649 39780 2659 40540
rect 2699 39780 2709 40540
rect 2649 39760 2709 39780
rect 2759 40540 2819 40620
rect 2759 39780 2769 40540
rect 2809 39780 2819 40540
rect 2869 40770 2929 40790
rect 2869 40730 2879 40770
rect 2919 40730 2929 40770
rect 2869 40530 2929 40730
rect 3089 40780 3149 40790
rect 3089 40740 3099 40780
rect 3139 40740 3149 40780
rect 2989 40660 3049 40680
rect 2989 40620 2999 40660
rect 3039 40620 3049 40660
rect 2989 40600 3049 40620
rect 2869 40490 2879 40530
rect 2919 40490 2929 40530
rect 2869 40470 2929 40490
rect 2979 40540 3039 40560
rect 2759 39760 2819 39780
rect 2979 39780 2989 40540
rect 3029 39780 3039 40540
rect 2649 39570 2699 39760
rect 2749 39690 2809 39710
rect 2749 39650 2759 39690
rect 2799 39650 2809 39690
rect 2749 39630 2809 39650
rect 2979 39570 3039 39780
rect 3089 40540 3149 40740
rect 4409 40780 4469 40790
rect 4409 40740 4419 40780
rect 4459 40740 4469 40780
rect 4409 40680 4469 40740
rect 4649 40680 4709 41080
rect 4759 41790 4819 41810
rect 4759 41080 4769 41790
rect 4809 41080 4819 41790
rect 4759 41060 4819 41080
rect 4869 41790 4929 41810
rect 4869 41080 4879 41790
rect 4919 41080 4929 41790
rect 4869 41060 4929 41080
rect 4979 41790 5039 41810
rect 4979 41080 4989 41790
rect 5029 41080 5039 41790
rect 4979 41060 5039 41080
rect 5089 41790 5149 41810
rect 5089 41080 5099 41790
rect 5139 41080 5149 41790
rect 5089 41060 5149 41080
rect 5199 41790 5259 41810
rect 5199 41080 5209 41790
rect 5249 41080 5259 41790
rect 5199 41060 5259 41080
rect 5309 41790 5369 41810
rect 5309 41080 5319 41790
rect 5359 41080 5369 41790
rect 5309 41060 5369 41080
rect 5419 41790 5479 41810
rect 5419 41080 5429 41790
rect 5469 41080 5479 41790
rect 5949 41360 5959 41820
rect 5999 41360 6009 41820
rect 5949 41340 6009 41360
rect 6059 41820 6119 41840
rect 6059 41360 6069 41820
rect 6109 41360 6119 41820
rect 5959 41280 6019 41300
rect 5959 41240 5969 41280
rect 6009 41240 6019 41280
rect 5959 41220 6019 41240
rect 6059 41280 6119 41360
rect 6179 41820 6239 41840
rect 6179 41360 6189 41820
rect 6229 41360 6239 41820
rect 6179 41340 6239 41360
rect 6289 41820 6349 41900
rect 6289 41360 6299 41820
rect 6339 41360 6349 41820
rect 6289 41340 6349 41360
rect 6399 41820 6459 41840
rect 6399 41360 6409 41820
rect 6449 41360 6459 41820
rect 6059 41240 6069 41280
rect 6109 41240 6119 41280
rect 5419 41060 5479 41080
rect 5949 41160 6009 41180
rect 5949 41000 5959 41160
rect 5999 41000 6009 41160
rect 5349 40980 5409 41000
rect 5349 40940 5359 40980
rect 5399 40940 5409 40980
rect 5349 40680 5409 40940
rect 5949 40920 6009 41000
rect 6059 41160 6119 41240
rect 6189 41280 6249 41300
rect 6189 41240 6199 41280
rect 6239 41240 6249 41280
rect 6189 41220 6249 41240
rect 6399 41280 6459 41360
rect 6519 41820 6579 41840
rect 6519 41360 6529 41820
rect 6569 41360 6579 41820
rect 6519 41340 6579 41360
rect 6629 41820 6689 41900
rect 6629 41360 6639 41820
rect 6679 41360 6689 41820
rect 6629 41340 6689 41360
rect 6739 41820 6799 41840
rect 6739 41360 6749 41820
rect 6789 41360 6799 41820
rect 6739 41340 6799 41360
rect 6849 41820 6909 41900
rect 6849 41360 6859 41820
rect 6899 41360 6909 41820
rect 6849 41340 6909 41360
rect 6959 41820 7019 41840
rect 6959 41360 6969 41820
rect 7009 41360 7019 41820
rect 6399 41240 6409 41280
rect 6449 41240 6459 41280
rect 6059 41000 6069 41160
rect 6109 41000 6119 41160
rect 6059 40980 6119 41000
rect 6179 41160 6239 41180
rect 6179 41000 6189 41160
rect 6229 41000 6239 41160
rect 6179 40980 6239 41000
rect 6289 41160 6349 41180
rect 6289 41000 6299 41160
rect 6339 41000 6349 41160
rect 6289 40920 6349 41000
rect 6399 41160 6459 41240
rect 6529 41280 6589 41300
rect 6529 41240 6539 41280
rect 6579 41240 6589 41280
rect 6529 41220 6589 41240
rect 6959 41280 7019 41360
rect 7079 41820 7139 41840
rect 7079 41360 7089 41820
rect 7129 41360 7139 41820
rect 7079 41340 7139 41360
rect 7189 41820 7249 41900
rect 7189 41360 7199 41820
rect 7239 41360 7249 41820
rect 7189 41340 7249 41360
rect 7299 41820 7359 41840
rect 7299 41360 7309 41820
rect 7349 41360 7359 41820
rect 7299 41340 7359 41360
rect 7409 41820 7469 41900
rect 7409 41360 7419 41820
rect 7459 41360 7469 41820
rect 7409 41340 7469 41360
rect 7519 41820 7579 41840
rect 7519 41360 7529 41820
rect 7569 41360 7579 41820
rect 7519 41340 7579 41360
rect 7629 41820 7689 41900
rect 7629 41360 7639 41820
rect 7679 41360 7689 41820
rect 7629 41340 7689 41360
rect 7739 41820 7799 41840
rect 7739 41360 7749 41820
rect 7789 41360 7799 41820
rect 7739 41340 7799 41360
rect 7849 41820 7909 41900
rect 7849 41360 7859 41820
rect 7899 41360 7909 41820
rect 7849 41340 7909 41360
rect 7959 41820 8019 41840
rect 7959 41360 7969 41820
rect 8009 41360 8019 41820
rect 6959 41240 6969 41280
rect 7009 41240 7019 41280
rect 6399 41000 6409 41160
rect 6449 41000 6459 41160
rect 6399 40980 6459 41000
rect 6519 41160 6579 41180
rect 6519 41000 6529 41160
rect 6569 41000 6579 41160
rect 6519 40980 6579 41000
rect 6629 41160 6689 41180
rect 6629 41000 6639 41160
rect 6679 41000 6689 41160
rect 6629 40920 6689 41000
rect 6739 41160 6799 41180
rect 6739 41000 6749 41160
rect 6789 41000 6799 41160
rect 6739 40980 6799 41000
rect 6849 41160 6909 41180
rect 6849 41000 6859 41160
rect 6899 41000 6909 41160
rect 6849 40920 6909 41000
rect 6959 41160 7019 41240
rect 7089 41280 7149 41300
rect 7089 41240 7099 41280
rect 7139 41240 7149 41280
rect 7089 41220 7149 41240
rect 7959 41280 8019 41360
rect 8139 41820 8199 41840
rect 8139 41360 8149 41820
rect 8189 41360 8199 41820
rect 8139 41340 8199 41360
rect 8249 41820 8309 41900
rect 8249 41360 8259 41820
rect 8299 41360 8309 41820
rect 8249 41340 8309 41360
rect 8359 41820 8419 41840
rect 8359 41360 8369 41820
rect 8409 41360 8419 41820
rect 8359 41340 8419 41360
rect 8469 41820 8529 41900
rect 8469 41360 8479 41820
rect 8519 41360 8529 41820
rect 8469 41340 8529 41360
rect 8579 41820 8639 41840
rect 8579 41360 8589 41820
rect 8629 41360 8639 41820
rect 8579 41340 8639 41360
rect 8689 41820 8749 41900
rect 8689 41360 8699 41820
rect 8739 41360 8749 41820
rect 8689 41340 8749 41360
rect 8799 41820 8859 41840
rect 8799 41360 8809 41820
rect 8849 41360 8859 41820
rect 8799 41340 8859 41360
rect 8909 41820 8969 41900
rect 8909 41360 8919 41820
rect 8959 41360 8969 41820
rect 8909 41340 8969 41360
rect 9019 41820 9079 41840
rect 9019 41360 9029 41820
rect 9069 41360 9079 41820
rect 9019 41340 9079 41360
rect 9129 41820 9189 41900
rect 9129 41360 9139 41820
rect 9179 41360 9189 41820
rect 9129 41340 9189 41360
rect 9239 41820 9299 41840
rect 9239 41360 9249 41820
rect 9289 41360 9299 41820
rect 9239 41340 9299 41360
rect 9349 41820 9409 41900
rect 9349 41360 9359 41820
rect 9399 41360 9409 41820
rect 9349 41340 9409 41360
rect 9459 41820 9519 41840
rect 9459 41360 9469 41820
rect 9509 41360 9519 41820
rect 9459 41340 9519 41360
rect 9569 41820 9629 41900
rect 9569 41360 9579 41820
rect 9619 41360 9629 41820
rect 9569 41340 9629 41360
rect 9679 41820 9739 41840
rect 9679 41360 9689 41820
rect 9729 41360 9739 41820
rect 9679 41340 9739 41360
rect 9789 41820 9849 41900
rect 21720 41860 21780 41900
rect 22580 41910 22940 41930
rect 23110 41970 23330 41990
rect 23110 41930 23120 41970
rect 23160 41930 23330 41970
rect 9789 41360 9799 41820
rect 9839 41360 9849 41820
rect 9789 41340 9849 41360
rect 9899 41820 9959 41840
rect 9899 41360 9909 41820
rect 9949 41360 9959 41820
rect 21720 41700 21730 41860
rect 21770 41700 21780 41860
rect 21720 41680 21780 41700
rect 21830 41860 21890 41880
rect 21830 41700 21840 41860
rect 21880 41700 21890 41860
rect 22580 41810 22630 41910
rect 22570 41800 22650 41810
rect 22570 41760 22590 41800
rect 22630 41760 22650 41800
rect 22570 41750 22650 41760
rect 7959 41240 7969 41280
rect 8009 41240 8019 41280
rect 6959 41000 6969 41160
rect 7009 41000 7019 41160
rect 6959 40980 7019 41000
rect 7079 41160 7139 41180
rect 7079 41000 7089 41160
rect 7129 41000 7139 41160
rect 7079 40980 7139 41000
rect 7189 41160 7249 41180
rect 7189 41000 7199 41160
rect 7239 41000 7249 41160
rect 7189 40920 7249 41000
rect 7299 41160 7359 41180
rect 7299 41000 7309 41160
rect 7349 41000 7359 41160
rect 7299 40980 7359 41000
rect 7409 41160 7469 41180
rect 7409 41000 7419 41160
rect 7459 41000 7469 41160
rect 7409 40920 7469 41000
rect 7519 41160 7579 41180
rect 7519 41000 7529 41160
rect 7569 41000 7579 41160
rect 7519 40980 7579 41000
rect 7629 41160 7689 41180
rect 7629 41000 7639 41160
rect 7679 41000 7689 41160
rect 7629 40920 7689 41000
rect 7739 41160 7799 41180
rect 7739 41000 7749 41160
rect 7789 41000 7799 41160
rect 7739 40980 7799 41000
rect 7849 41160 7909 41180
rect 7849 41000 7859 41160
rect 7899 41000 7909 41160
rect 7849 40920 7909 41000
rect 7959 41160 8019 41240
rect 8149 41280 8209 41300
rect 8149 41240 8159 41280
rect 8199 41240 8209 41280
rect 8149 41220 8209 41240
rect 9899 41290 9959 41360
rect 9899 41280 10029 41290
rect 9899 41230 9959 41280
rect 10009 41230 10029 41280
rect 9899 41220 10029 41230
rect 7959 41000 7969 41160
rect 8009 41000 8019 41160
rect 7959 40980 8019 41000
rect 8139 41160 8199 41180
rect 8139 41000 8149 41160
rect 8189 41000 8199 41160
rect 8139 40980 8199 41000
rect 8249 41160 8309 41180
rect 8249 41000 8259 41160
rect 8299 41000 8309 41160
rect 8249 40920 8309 41000
rect 8359 41160 8419 41180
rect 8359 41000 8369 41160
rect 8409 41000 8419 41160
rect 8359 40980 8419 41000
rect 8469 41160 8529 41180
rect 8469 41000 8479 41160
rect 8519 41000 8529 41160
rect 8469 40920 8529 41000
rect 8579 41160 8639 41180
rect 8579 41000 8589 41160
rect 8629 41000 8639 41160
rect 8579 40980 8639 41000
rect 8689 41160 8749 41180
rect 8689 41000 8699 41160
rect 8739 41000 8749 41160
rect 8689 40920 8749 41000
rect 8799 41160 8859 41180
rect 8799 41000 8809 41160
rect 8849 41000 8859 41160
rect 8799 40980 8859 41000
rect 8909 41160 8969 41180
rect 8909 41000 8919 41160
rect 8959 41000 8969 41160
rect 8909 40920 8969 41000
rect 9019 41160 9079 41180
rect 9019 41000 9029 41160
rect 9069 41000 9079 41160
rect 9019 40980 9079 41000
rect 9129 41160 9189 41180
rect 9129 41000 9139 41160
rect 9179 41000 9189 41160
rect 9129 40920 9189 41000
rect 9239 41160 9299 41180
rect 9239 41000 9249 41160
rect 9289 41000 9299 41160
rect 9239 40980 9299 41000
rect 9349 41160 9409 41180
rect 9349 41000 9359 41160
rect 9399 41000 9409 41160
rect 9349 40920 9409 41000
rect 9459 41160 9519 41180
rect 9459 41000 9469 41160
rect 9509 41000 9519 41160
rect 9459 40980 9519 41000
rect 9569 41160 9629 41180
rect 9569 41000 9579 41160
rect 9619 41000 9629 41160
rect 9569 40920 9629 41000
rect 9679 41160 9739 41180
rect 9679 41000 9689 41160
rect 9729 41000 9739 41160
rect 9679 40980 9739 41000
rect 9789 41160 9849 41180
rect 9789 41000 9799 41160
rect 9839 41000 9849 41160
rect 9789 40920 9849 41000
rect 9899 41160 9959 41220
rect 21830 41180 21890 41700
rect 22580 41690 22640 41710
rect 22580 41530 22590 41690
rect 22630 41530 22640 41690
rect 22430 41330 22530 41350
rect 22580 41330 22640 41530
rect 22430 41270 22450 41330
rect 22510 41270 22640 41330
rect 22690 41690 22750 41710
rect 22690 41530 22700 41690
rect 22740 41530 22750 41690
rect 22690 41310 22750 41530
rect 22880 41690 22940 41910
rect 22980 41910 23060 41920
rect 23110 41910 23330 41930
rect 22980 41870 23000 41910
rect 23040 41870 23150 41910
rect 22980 41860 23060 41870
rect 23110 41810 23150 41870
rect 23280 41860 23330 41910
rect 23380 42080 23440 42100
rect 23380 41920 23390 42080
rect 23430 41920 23440 42080
rect 23380 41860 23440 41920
rect 23280 41810 23440 41860
rect 23490 42080 23550 42100
rect 23490 41920 23500 42080
rect 23540 41920 23550 42080
rect 23490 41870 23550 41920
rect 23620 41870 23740 41890
rect 23490 41810 23640 41870
rect 23720 41810 23740 41870
rect 23090 41800 23170 41810
rect 23090 41760 23110 41800
rect 23150 41760 23170 41800
rect 23090 41750 23170 41760
rect 22880 41530 22890 41690
rect 22930 41530 22940 41690
rect 22880 41510 22940 41530
rect 22990 41690 23050 41710
rect 22990 41530 23000 41690
rect 23040 41530 23050 41690
rect 22990 41310 23050 41530
rect 22430 41250 22530 41270
rect 22690 41260 23050 41310
rect 23100 41690 23160 41710
rect 23100 41530 23110 41690
rect 23150 41530 23160 41690
rect 23100 41180 23160 41530
rect 23280 41290 23330 41810
rect 23490 41770 23550 41810
rect 23620 41790 23740 41810
rect 23480 41760 23560 41770
rect 23480 41720 23500 41760
rect 23540 41720 23560 41760
rect 23480 41710 23560 41720
rect 23800 41690 23880 41710
rect 23800 41670 23810 41690
rect 23380 41630 23810 41670
rect 23870 41630 23880 41690
rect 23380 41610 23880 41630
rect 23380 41550 23440 41610
rect 23380 41390 23390 41550
rect 23430 41390 23440 41550
rect 23380 41370 23440 41390
rect 23490 41550 23550 41570
rect 23490 41390 23500 41550
rect 23540 41390 23550 41550
rect 23490 41290 23550 41390
rect 23280 41230 23550 41290
rect 9899 41000 9909 41160
rect 9949 41000 9959 41160
rect 21590 41160 23630 41180
rect 21590 41090 21620 41160
rect 21680 41090 21720 41160
rect 21780 41090 21830 41160
rect 21890 41090 21930 41160
rect 21990 41090 22030 41160
rect 22090 41090 22130 41160
rect 22190 41090 22230 41160
rect 22290 41090 22330 41160
rect 22390 41090 22430 41160
rect 22490 41090 22530 41160
rect 22590 41090 22630 41160
rect 22690 41090 22730 41160
rect 22790 41090 22830 41160
rect 22890 41090 22930 41160
rect 22990 41090 23030 41160
rect 23090 41090 23130 41160
rect 23190 41090 23230 41160
rect 23290 41090 23330 41160
rect 23390 41090 23430 41160
rect 23490 41090 23530 41160
rect 23590 41090 23630 41160
rect 21590 41080 23630 41090
rect 9899 40980 9959 41000
rect 5949 40910 9979 40920
rect 5949 40850 6009 40910
rect 6070 40850 9979 40910
rect 5949 40840 9979 40850
rect 5449 40780 5519 40790
rect 5449 40740 5459 40780
rect 5499 40740 5519 40780
rect 5449 40730 5519 40740
rect 3089 39780 3099 40540
rect 3139 39780 3149 40540
rect 3260 40670 4469 40680
rect 3260 40610 3320 40670
rect 3380 40610 3430 40670
rect 3490 40610 3540 40670
rect 3600 40610 3650 40670
rect 3710 40610 3760 40670
rect 3820 40610 3870 40670
rect 3930 40610 3980 40670
rect 4040 40610 4090 40670
rect 4150 40610 4469 40670
rect 3260 40600 4469 40610
rect 3260 40530 3319 40600
rect 3260 40510 3320 40530
rect 3260 39800 3269 40510
rect 3309 39800 3320 40510
rect 3260 39780 3320 39800
rect 3369 40510 3430 40530
rect 3369 39800 3379 40510
rect 3419 39800 3430 40510
rect 3369 39780 3430 39800
rect 3479 40510 3540 40530
rect 3479 39800 3489 40510
rect 3529 39800 3540 40510
rect 3479 39780 3540 39800
rect 3589 40510 3650 40530
rect 3589 39800 3599 40510
rect 3639 39800 3650 40510
rect 3589 39780 3650 39800
rect 3699 40510 3760 40530
rect 3699 39800 3709 40510
rect 3749 39800 3760 40510
rect 3699 39780 3760 39800
rect 3809 40510 3870 40530
rect 3809 39800 3819 40510
rect 3859 39800 3870 40510
rect 3809 39780 3870 39800
rect 3919 40510 3980 40530
rect 3919 39800 3929 40510
rect 3969 39800 3980 40510
rect 3919 39780 3980 39800
rect 4029 40510 4090 40530
rect 4029 39800 4039 40510
rect 4079 39800 4090 40510
rect 4029 39780 4090 39800
rect 4139 40510 4200 40530
rect 4139 39800 4149 40510
rect 4189 39800 4200 40510
rect 4139 39780 4200 39800
rect 3089 39760 3149 39780
rect 3329 39700 3389 39720
rect 3329 39660 3339 39700
rect 3379 39660 3389 39700
rect 3329 39640 3389 39660
rect 4029 39570 4089 39780
rect 4409 39690 4469 40600
rect 4539 40660 5429 40680
rect 4539 40620 4659 40660
rect 5399 40620 5429 40660
rect 4539 40600 5429 40620
rect 6349 40650 9969 40660
rect 4539 40510 4599 40600
rect 6349 40590 6409 40650
rect 6469 40590 6519 40650
rect 6579 40590 6629 40650
rect 6689 40590 6739 40650
rect 6799 40590 6849 40650
rect 6909 40590 6959 40650
rect 7019 40590 7069 40650
rect 7129 40590 7179 40650
rect 7239 40590 7289 40650
rect 7349 40590 7399 40650
rect 7459 40590 7509 40650
rect 7569 40590 7619 40650
rect 7679 40590 7729 40650
rect 7789 40590 7839 40650
rect 7899 40590 7949 40650
rect 8009 40590 8059 40650
rect 8119 40590 8169 40650
rect 8229 40590 8279 40650
rect 8339 40590 8389 40650
rect 8449 40590 8499 40650
rect 8559 40590 8609 40650
rect 8669 40590 8719 40650
rect 8779 40590 8829 40650
rect 8889 40590 8939 40650
rect 8999 40590 9049 40650
rect 9109 40590 9159 40650
rect 9219 40590 9269 40650
rect 9329 40590 9379 40650
rect 9439 40590 9489 40650
rect 9549 40590 9599 40650
rect 9659 40590 9709 40650
rect 9769 40590 9819 40650
rect 9879 40590 9969 40650
rect 6349 40580 9969 40590
rect 4539 39800 4549 40510
rect 4589 39800 4599 40510
rect 4539 39780 4599 39800
rect 4649 40510 4709 40530
rect 4649 39800 4659 40510
rect 4699 39800 4709 40510
rect 4649 39690 4709 39800
rect 4759 40510 4819 40530
rect 4759 39800 4769 40510
rect 4809 39800 4819 40510
rect 4759 39780 4819 39800
rect 4869 40510 4929 40530
rect 4869 39800 4879 40510
rect 4919 39800 4929 40510
rect 4869 39780 4929 39800
rect 4979 40510 5039 40530
rect 4979 39800 4989 40510
rect 5029 39800 5039 40510
rect 4979 39780 5039 39800
rect 5089 40510 5149 40530
rect 5089 39800 5099 40510
rect 5139 39800 5149 40510
rect 5089 39780 5149 39800
rect 5199 40510 5259 40530
rect 5199 39800 5209 40510
rect 5249 39800 5259 40510
rect 5199 39780 5259 39800
rect 5309 40510 5369 40530
rect 5309 39800 5319 40510
rect 5359 39800 5369 40510
rect 5309 39780 5369 39800
rect 5419 40510 5479 40530
rect 5419 39800 5429 40510
rect 5469 39800 5479 40510
rect 6349 40500 6409 40520
rect 6349 40040 6359 40500
rect 6399 40040 6409 40500
rect 6349 40020 6409 40040
rect 6459 40500 6519 40580
rect 6459 40040 6469 40500
rect 6509 40040 6519 40500
rect 6459 40020 6519 40040
rect 6569 40500 6629 40520
rect 6569 40040 6579 40500
rect 6619 40040 6629 40500
rect 6569 40020 6629 40040
rect 6679 40500 6739 40580
rect 6679 40040 6689 40500
rect 6729 40040 6739 40500
rect 6679 40020 6739 40040
rect 6789 40500 6849 40520
rect 6789 40040 6799 40500
rect 6839 40040 6849 40500
rect 6789 40020 6849 40040
rect 6899 40500 6959 40580
rect 6899 40040 6909 40500
rect 6949 40040 6959 40500
rect 6899 40020 6959 40040
rect 7009 40500 7069 40520
rect 7009 40040 7019 40500
rect 7059 40040 7069 40500
rect 7009 40020 7069 40040
rect 7119 40500 7179 40580
rect 7119 40040 7129 40500
rect 7169 40040 7179 40500
rect 7119 40020 7179 40040
rect 7229 40500 7289 40520
rect 7229 40040 7239 40500
rect 7279 40040 7289 40500
rect 7229 40020 7289 40040
rect 7339 40500 7399 40580
rect 7339 40040 7349 40500
rect 7389 40040 7399 40500
rect 7339 40020 7399 40040
rect 7449 40500 7509 40520
rect 7449 40040 7459 40500
rect 7499 40040 7509 40500
rect 7449 40020 7509 40040
rect 7559 40500 7619 40580
rect 7559 40040 7569 40500
rect 7609 40040 7619 40500
rect 7559 40020 7619 40040
rect 7669 40500 7729 40520
rect 7669 40040 7679 40500
rect 7719 40040 7729 40500
rect 7669 40020 7729 40040
rect 7779 40500 7839 40580
rect 7779 40040 7789 40500
rect 7829 40040 7839 40500
rect 7779 40020 7839 40040
rect 7889 40500 7949 40520
rect 7889 40040 7899 40500
rect 7939 40040 7949 40500
rect 7889 40020 7949 40040
rect 7999 40500 8059 40580
rect 7999 40040 8009 40500
rect 8049 40040 8059 40500
rect 7999 40020 8059 40040
rect 8109 40500 8169 40520
rect 8109 40040 8119 40500
rect 8159 40040 8169 40500
rect 8109 40020 8169 40040
rect 8219 40500 8279 40580
rect 8219 40040 8229 40500
rect 8269 40040 8279 40500
rect 8219 40020 8279 40040
rect 8329 40500 8389 40520
rect 8329 40040 8339 40500
rect 8379 40040 8389 40500
rect 8329 40020 8389 40040
rect 8439 40500 8499 40580
rect 8439 40040 8449 40500
rect 8489 40040 8499 40500
rect 8439 40020 8499 40040
rect 8549 40500 8609 40520
rect 8549 40040 8559 40500
rect 8599 40040 8609 40500
rect 8549 40020 8609 40040
rect 8659 40500 8719 40580
rect 8659 40040 8669 40500
rect 8709 40040 8719 40500
rect 8659 40020 8719 40040
rect 8769 40500 8829 40520
rect 8769 40040 8779 40500
rect 8819 40040 8829 40500
rect 8769 40020 8829 40040
rect 8879 40500 8939 40580
rect 8879 40040 8889 40500
rect 8929 40040 8939 40500
rect 8879 40020 8939 40040
rect 8989 40500 9049 40520
rect 8989 40040 8999 40500
rect 9039 40040 9049 40500
rect 8989 40020 9049 40040
rect 9099 40500 9159 40580
rect 9099 40040 9109 40500
rect 9149 40040 9159 40500
rect 9099 40020 9159 40040
rect 9209 40500 9269 40520
rect 9209 40040 9219 40500
rect 9259 40040 9269 40500
rect 9209 40020 9269 40040
rect 9319 40500 9379 40580
rect 9319 40040 9329 40500
rect 9369 40040 9379 40500
rect 9319 40020 9379 40040
rect 9429 40500 9489 40520
rect 9429 40040 9439 40500
rect 9479 40040 9489 40500
rect 9429 40020 9489 40040
rect 9539 40500 9599 40580
rect 9539 40040 9549 40500
rect 9589 40040 9599 40500
rect 9539 40020 9599 40040
rect 9649 40500 9709 40520
rect 9649 40040 9659 40500
rect 9699 40040 9709 40500
rect 9649 40020 9709 40040
rect 9759 40500 9819 40580
rect 9759 40040 9769 40500
rect 9809 40040 9819 40500
rect 9759 40020 9819 40040
rect 9869 40500 9929 40520
rect 9869 40040 9879 40500
rect 9919 40040 9929 40500
rect 6349 39960 6419 39980
rect 6349 39920 6369 39960
rect 6409 39920 6419 39960
rect 6349 39900 6419 39920
rect 9869 39970 9929 40040
rect 9869 39960 9999 39970
rect 9869 39910 9929 39960
rect 9979 39910 9999 39960
rect 9869 39900 9999 39910
rect 5419 39780 5479 39800
rect 6349 39840 6409 39860
rect 4409 39650 4709 39690
rect 5349 39700 5409 39720
rect 5349 39660 5359 39700
rect 5399 39660 5409 39700
rect 6349 39680 6359 39840
rect 6399 39680 6409 39840
rect 6349 39660 6409 39680
rect 6459 39840 6519 39860
rect 6459 39680 6469 39840
rect 6509 39680 6519 39840
rect 5349 39640 5409 39660
rect 6459 39570 6519 39680
rect 6569 39840 6629 39860
rect 6569 39680 6579 39840
rect 6619 39680 6629 39840
rect 6569 39660 6629 39680
rect 6679 39840 6739 39860
rect 6679 39680 6689 39840
rect 6729 39680 6739 39840
rect 6679 39570 6739 39680
rect 6789 39840 6849 39860
rect 6789 39680 6799 39840
rect 6839 39680 6849 39840
rect 6789 39660 6849 39680
rect 6899 39840 6959 39860
rect 6899 39680 6909 39840
rect 6949 39680 6959 39840
rect 6899 39570 6959 39680
rect 7009 39840 7069 39860
rect 7009 39680 7019 39840
rect 7059 39680 7069 39840
rect 7009 39660 7069 39680
rect 7119 39840 7179 39860
rect 7119 39680 7129 39840
rect 7169 39680 7179 39840
rect 7119 39570 7179 39680
rect 7229 39840 7289 39860
rect 7229 39680 7239 39840
rect 7279 39680 7289 39840
rect 7229 39660 7289 39680
rect 7339 39840 7399 39860
rect 7339 39680 7349 39840
rect 7389 39680 7399 39840
rect 7339 39570 7399 39680
rect 7449 39840 7509 39860
rect 7449 39680 7459 39840
rect 7499 39680 7509 39840
rect 7449 39660 7509 39680
rect 7559 39840 7619 39860
rect 7559 39680 7569 39840
rect 7609 39680 7619 39840
rect 7559 39570 7619 39680
rect 7669 39840 7729 39860
rect 7669 39680 7679 39840
rect 7719 39680 7729 39840
rect 7669 39660 7729 39680
rect 7779 39840 7839 39860
rect 7779 39680 7789 39840
rect 7829 39680 7839 39840
rect 7779 39570 7839 39680
rect 7889 39840 7949 39860
rect 7889 39680 7899 39840
rect 7939 39680 7949 39840
rect 7889 39660 7949 39680
rect 7999 39840 8059 39860
rect 7999 39680 8009 39840
rect 8049 39680 8059 39840
rect 7999 39570 8059 39680
rect 8109 39840 8169 39860
rect 8109 39680 8119 39840
rect 8159 39680 8169 39840
rect 8109 39660 8169 39680
rect 8219 39840 8279 39860
rect 8219 39680 8229 39840
rect 8269 39680 8279 39840
rect 8219 39570 8279 39680
rect 8329 39840 8389 39860
rect 8329 39680 8339 39840
rect 8379 39680 8389 39840
rect 8329 39660 8389 39680
rect 8439 39840 8499 39860
rect 8439 39680 8449 39840
rect 8489 39680 8499 39840
rect 8439 39570 8499 39680
rect 8549 39840 8609 39860
rect 8549 39680 8559 39840
rect 8599 39680 8609 39840
rect 8549 39660 8609 39680
rect 8659 39840 8719 39860
rect 8659 39680 8669 39840
rect 8709 39680 8719 39840
rect 8659 39570 8719 39680
rect 8769 39840 8829 39860
rect 8769 39680 8779 39840
rect 8819 39680 8829 39840
rect 8769 39660 8829 39680
rect 8879 39840 8939 39860
rect 8879 39680 8889 39840
rect 8929 39680 8939 39840
rect 8879 39570 8939 39680
rect 8989 39840 9049 39860
rect 8989 39680 8999 39840
rect 9039 39680 9049 39840
rect 8989 39660 9049 39680
rect 9099 39840 9159 39860
rect 9099 39680 9109 39840
rect 9149 39680 9159 39840
rect 9099 39570 9159 39680
rect 9209 39840 9269 39860
rect 9209 39680 9219 39840
rect 9259 39680 9269 39840
rect 9209 39660 9269 39680
rect 9319 39840 9379 39860
rect 9319 39680 9329 39840
rect 9369 39680 9379 39840
rect 9319 39570 9379 39680
rect 9429 39840 9489 39860
rect 9429 39680 9439 39840
rect 9479 39680 9489 39840
rect 9429 39660 9489 39680
rect 9539 39840 9599 39860
rect 9539 39680 9549 39840
rect 9589 39680 9599 39840
rect 9539 39570 9599 39680
rect 9649 39840 9709 39860
rect 9649 39680 9659 39840
rect 9699 39680 9709 39840
rect 9649 39660 9709 39680
rect 9759 39840 9819 39860
rect 9759 39680 9769 39840
rect 9809 39680 9819 39840
rect 9759 39570 9819 39680
rect 9869 39840 9929 39900
rect 9869 39680 9879 39840
rect 9919 39680 9929 39840
rect 9869 39660 9929 39680
rect 2619 39560 9979 39570
rect 2619 39500 2649 39560
rect 2709 39500 2749 39560
rect 2809 39500 2849 39560
rect 2909 39500 2949 39560
rect 3009 39500 3049 39560
rect 3109 39500 3149 39560
rect 3209 39500 3249 39560
rect 3309 39500 3349 39560
rect 3409 39500 3449 39560
rect 3509 39500 3549 39560
rect 3609 39500 3649 39560
rect 3709 39500 3749 39560
rect 3809 39500 3849 39560
rect 3909 39500 3949 39560
rect 4009 39500 4049 39560
rect 4109 39500 4149 39560
rect 4209 39500 4249 39560
rect 4309 39500 4349 39560
rect 4409 39500 4449 39560
rect 4509 39500 4549 39560
rect 4609 39500 4649 39560
rect 4709 39500 4749 39560
rect 4809 39500 4849 39560
rect 4909 39500 4949 39560
rect 5009 39500 5049 39560
rect 5109 39500 5149 39560
rect 5209 39500 5249 39560
rect 5309 39500 6349 39560
rect 6409 39500 6449 39560
rect 6509 39500 6549 39560
rect 6609 39500 6649 39560
rect 6709 39500 6749 39560
rect 6809 39500 6849 39560
rect 6909 39500 6949 39560
rect 7009 39500 7049 39560
rect 7109 39500 7149 39560
rect 7209 39500 7249 39560
rect 7309 39500 7349 39560
rect 7409 39500 7479 39560
rect 7539 39500 7579 39560
rect 7639 39500 7679 39560
rect 7739 39500 7779 39560
rect 7839 39500 7879 39560
rect 7939 39500 7979 39560
rect 8039 39500 8079 39560
rect 8139 39500 8179 39560
rect 8239 39500 8279 39560
rect 8339 39500 8379 39560
rect 8439 39500 8479 39560
rect 8539 39500 8629 39560
rect 8689 39500 8729 39560
rect 8789 39500 8829 39560
rect 8889 39500 8929 39560
rect 8989 39500 9029 39560
rect 9089 39500 9129 39560
rect 9189 39500 9229 39560
rect 9289 39500 9329 39560
rect 9389 39500 9429 39560
rect 9489 39500 9529 39560
rect 9589 39500 9629 39560
rect 9689 39500 9739 39560
rect 9799 39500 9839 39560
rect 9899 39500 9979 39560
rect 2619 39490 9979 39500
rect 3770 37180 6200 37190
rect 3770 37120 3810 37180
rect 3870 37120 3910 37180
rect 3970 37120 4010 37180
rect 4070 37120 4110 37180
rect 4170 37120 4210 37180
rect 4270 37120 4310 37180
rect 4370 37120 4410 37180
rect 4470 37120 4510 37180
rect 4570 37120 4610 37180
rect 4670 37120 4710 37180
rect 4770 37120 4810 37180
rect 4870 37120 4910 37180
rect 4970 37120 5010 37180
rect 5070 37120 5110 37180
rect 5170 37120 5210 37180
rect 5270 37120 5310 37180
rect 5370 37120 5410 37180
rect 5470 37120 5510 37180
rect 5570 37120 5610 37180
rect 5670 37120 5710 37180
rect 5770 37120 5810 37180
rect 5870 37120 5910 37180
rect 5970 37120 6010 37180
rect 6070 37120 6110 37180
rect 6170 37120 6200 37180
rect 3770 37110 6200 37120
rect 3770 37030 3830 37110
rect 3770 36270 3780 37030
rect 3820 36270 3830 37030
rect 3770 36250 3830 36270
rect 3880 37030 3940 37050
rect 3880 36270 3890 37030
rect 3930 36270 3940 37030
rect 3880 36250 3940 36270
rect 3990 37030 4050 37050
rect 3990 36270 4000 37030
rect 4040 36270 4050 37030
rect 3990 36250 4050 36270
rect 4100 37030 4160 37050
rect 4100 36270 4110 37030
rect 4150 36270 4160 37030
rect 4100 36250 4160 36270
rect 4210 37030 4270 37050
rect 4210 36270 4220 37030
rect 4260 36270 4270 37030
rect 4210 36250 4270 36270
rect 4320 37030 4380 37050
rect 4320 36270 4330 37030
rect 4370 36270 4380 37030
rect 4320 36250 4380 36270
rect 4500 37030 4560 37050
rect 4500 36270 4510 37030
rect 4550 36270 4560 37030
rect 4500 36250 4560 36270
rect 4690 37030 4750 37050
rect 4690 36270 4700 37030
rect 4740 36270 4750 37030
rect 4690 36250 4750 36270
rect 4800 37030 4860 37050
rect 4800 36270 4810 37030
rect 4850 36270 4860 37030
rect 4800 36250 4860 36270
rect 4910 37030 4970 37050
rect 4910 36270 4920 37030
rect 4960 36270 4970 37030
rect 4910 36250 4970 36270
rect 5020 37030 5080 37050
rect 5020 36270 5030 37030
rect 5070 36270 5080 37030
rect 5020 36250 5080 36270
rect 5130 37030 5190 37050
rect 5130 36270 5140 37030
rect 5180 36270 5190 37030
rect 5130 36250 5190 36270
rect 5240 37030 5300 37050
rect 5240 36270 5250 37030
rect 5290 36270 5300 37030
rect 5460 37030 5520 37050
rect 5460 36670 5470 37030
rect 5510 36670 5520 37030
rect 5460 36650 5520 36670
rect 5570 37030 5630 37110
rect 5570 36670 5580 37030
rect 5620 36670 5630 37030
rect 5570 36650 5630 36670
rect 5680 37030 5740 37050
rect 5680 36670 5690 37030
rect 5730 36670 5740 37030
rect 5680 36650 5740 36670
rect 5790 37030 5850 37110
rect 5790 36670 5800 37030
rect 5840 36670 5850 37030
rect 5790 36650 5850 36670
rect 5900 37030 5960 37050
rect 5900 36670 5910 37030
rect 5950 36670 5960 37030
rect 5900 36650 5960 36670
rect 6010 37030 6070 37110
rect 6010 36670 6020 37030
rect 6060 36670 6070 37030
rect 6010 36650 6070 36670
rect 6120 37030 6180 37050
rect 6120 36670 6130 37030
rect 6170 36670 6180 37030
rect 3730 34990 3840 35010
rect 3730 34940 3760 34990
rect 3810 34940 3840 34990
rect 3730 34920 3840 34940
rect 4530 35000 4650 35010
rect 4530 34930 4560 35000
rect 4620 34930 4650 35000
rect 4530 34920 4650 34930
rect 5240 34890 5300 36270
rect 5240 34870 5530 34890
rect 3770 34820 5310 34870
rect 5360 34820 5420 34870
rect 5470 34820 5530 34870
rect 3770 34800 5530 34820
rect 6120 34870 6180 36670
rect 6340 36720 10880 36730
rect 6340 36660 6380 36720
rect 6440 36660 6480 36720
rect 6540 36660 6580 36720
rect 6640 36660 6680 36720
rect 6740 36660 6780 36720
rect 6840 36660 6880 36720
rect 6940 36660 6980 36720
rect 7040 36660 7080 36720
rect 7140 36660 7180 36720
rect 7240 36660 7280 36720
rect 7340 36660 7380 36720
rect 7440 36660 7480 36720
rect 7540 36660 7580 36720
rect 7640 36660 7680 36720
rect 7740 36660 7780 36720
rect 7840 36660 7880 36720
rect 7940 36660 7980 36720
rect 8040 36660 8080 36720
rect 8140 36660 8180 36720
rect 8240 36660 8280 36720
rect 8340 36660 8380 36720
rect 8440 36660 8480 36720
rect 8540 36660 8580 36720
rect 8640 36660 8680 36720
rect 8740 36660 8780 36720
rect 8840 36660 8880 36720
rect 8940 36660 8980 36720
rect 9040 36660 9080 36720
rect 9140 36660 9180 36720
rect 9240 36660 9280 36720
rect 9340 36660 9380 36720
rect 9440 36660 9480 36720
rect 9540 36660 9580 36720
rect 9640 36660 9680 36720
rect 9740 36660 9780 36720
rect 9840 36660 9880 36720
rect 9940 36660 9980 36720
rect 10040 36660 10080 36720
rect 10140 36660 10180 36720
rect 10240 36660 10280 36720
rect 10340 36660 10380 36720
rect 10440 36660 10480 36720
rect 10540 36660 10580 36720
rect 10640 36660 10680 36720
rect 10740 36660 10780 36720
rect 10840 36660 10880 36720
rect 6340 36650 10880 36660
rect 6340 36570 6400 36650
rect 6340 36410 6350 36570
rect 6390 36410 6400 36570
rect 6340 36390 6400 36410
rect 6450 36570 6510 36590
rect 6450 36410 6460 36570
rect 6500 36410 6510 36570
rect 6120 34860 6260 34870
rect 6450 34860 6510 36410
rect 6560 36570 6620 36650
rect 6560 36410 6570 36570
rect 6610 36410 6620 36570
rect 6560 36390 6620 36410
rect 6810 36570 6870 36650
rect 6810 36210 6820 36570
rect 6860 36210 6870 36570
rect 6810 36190 6870 36210
rect 7070 36570 7130 36590
rect 7070 36210 7080 36570
rect 7120 36210 7130 36570
rect 7300 36570 7360 36650
rect 7300 36410 7310 36570
rect 7350 36410 7360 36570
rect 7300 36390 7360 36410
rect 7410 36570 7470 36590
rect 7410 36410 7420 36570
rect 7460 36410 7470 36570
rect 6710 34860 6770 34870
rect 6120 34810 6190 34860
rect 6240 34810 6260 34860
rect 6120 34800 6260 34810
rect 6320 34850 6410 34860
rect 6320 34810 6340 34850
rect 6380 34810 6410 34850
rect 6320 34800 6410 34810
rect 6450 34850 6770 34860
rect 7070 34850 7130 36210
rect 7410 34850 7470 36410
rect 7520 36570 7580 36650
rect 7520 36410 7530 36570
rect 7570 36410 7580 36570
rect 7520 36390 7580 36410
rect 7680 36570 7740 36650
rect 7680 36410 7690 36570
rect 7730 36410 7740 36570
rect 7680 36390 7740 36410
rect 7790 36570 7850 36590
rect 7790 36410 7800 36570
rect 7840 36410 7850 36570
rect 7790 34850 7850 36410
rect 7900 36570 7960 36650
rect 7900 36410 7910 36570
rect 7950 36410 7960 36570
rect 7900 36390 7960 36410
rect 8060 36570 8120 36650
rect 8060 36410 8070 36570
rect 8110 36410 8120 36570
rect 8060 36390 8120 36410
rect 8170 36570 8230 36590
rect 8170 36410 8180 36570
rect 8220 36410 8230 36570
rect 8170 34850 8230 36410
rect 8280 36570 8340 36650
rect 8280 36410 8290 36570
rect 8330 36410 8340 36570
rect 8280 36390 8340 36410
rect 8440 36570 8500 36650
rect 8440 36410 8450 36570
rect 8490 36410 8500 36570
rect 8440 36390 8500 36410
rect 8550 36570 8610 36590
rect 8550 36410 8560 36570
rect 8600 36410 8610 36570
rect 8550 34850 8610 36410
rect 8660 36570 8720 36650
rect 8660 36410 8670 36570
rect 8710 36410 8720 36570
rect 8660 36390 8720 36410
rect 8890 36570 8950 36650
rect 8890 36210 8900 36570
rect 8940 36210 8950 36570
rect 8890 36190 8950 36210
rect 9150 36570 9210 36590
rect 9150 36210 9160 36570
rect 9200 36210 9210 36570
rect 9380 36570 9440 36650
rect 9380 36410 9390 36570
rect 9430 36410 9440 36570
rect 9380 36390 9440 36410
rect 9490 36570 9550 36590
rect 9490 36410 9500 36570
rect 9540 36410 9550 36570
rect 8660 35460 8780 35500
rect 8660 35370 8680 35460
rect 8760 35370 8780 35460
rect 8660 35330 8780 35370
rect 8680 34850 8750 35330
rect 9050 34950 9110 34970
rect 9050 34910 9060 34950
rect 9100 34910 9110 34950
rect 9050 34890 9110 34910
rect 8790 34850 8850 34860
rect 9150 34850 9210 36210
rect 9490 34850 9550 36410
rect 9600 36570 9660 36650
rect 9600 36410 9610 36570
rect 9650 36410 9660 36570
rect 9600 36390 9660 36410
rect 9760 36570 9820 36650
rect 9760 36410 9770 36570
rect 9810 36410 9820 36570
rect 9760 36390 9820 36410
rect 9870 36570 9930 36590
rect 9870 36410 9880 36570
rect 9920 36410 9930 36570
rect 9870 34850 9930 36410
rect 9980 36570 10040 36650
rect 9980 36410 9990 36570
rect 10030 36410 10040 36570
rect 9980 36390 10040 36410
rect 10140 36570 10200 36650
rect 10140 36410 10150 36570
rect 10190 36410 10200 36570
rect 10140 36390 10200 36410
rect 10250 36570 10310 36590
rect 10250 36410 10260 36570
rect 10300 36410 10310 36570
rect 10250 34850 10310 36410
rect 10360 36570 10420 36650
rect 10360 36410 10370 36570
rect 10410 36410 10420 36570
rect 10360 36390 10420 36410
rect 10520 36570 10580 36650
rect 10520 36410 10530 36570
rect 10570 36410 10580 36570
rect 10520 36390 10580 36410
rect 10630 36570 10690 36590
rect 10630 36410 10640 36570
rect 10680 36410 10690 36570
rect 10630 34850 10690 36410
rect 10740 36570 10800 36650
rect 10740 36410 10750 36570
rect 10790 36410 10800 36570
rect 10740 36390 10800 36410
rect 15180 36340 24910 36350
rect 15180 36270 15220 36340
rect 15280 36270 15320 36340
rect 15380 36270 15420 36340
rect 15480 36270 15520 36340
rect 15580 36270 15620 36340
rect 15680 36270 15720 36340
rect 15780 36270 15820 36340
rect 15880 36270 15920 36340
rect 15980 36270 16020 36340
rect 16080 36270 16120 36340
rect 16180 36270 16220 36340
rect 16280 36270 16320 36340
rect 16380 36270 16420 36340
rect 16480 36270 16520 36340
rect 16580 36270 16620 36340
rect 16680 36270 16720 36340
rect 16780 36270 16820 36340
rect 16880 36270 16920 36340
rect 16980 36270 17020 36340
rect 17080 36270 17120 36340
rect 17180 36270 17220 36340
rect 17280 36270 17320 36340
rect 17380 36270 17420 36340
rect 17480 36270 17520 36340
rect 17580 36270 17620 36340
rect 17680 36270 17720 36340
rect 17780 36270 17820 36340
rect 17880 36270 17920 36340
rect 17980 36270 18020 36340
rect 18080 36270 18120 36340
rect 18180 36270 18220 36340
rect 18280 36270 18320 36340
rect 18380 36270 18420 36340
rect 18480 36270 18520 36340
rect 18580 36270 18620 36340
rect 18680 36270 18720 36340
rect 18780 36270 18820 36340
rect 18880 36270 18920 36340
rect 18980 36270 19020 36340
rect 19080 36270 19120 36340
rect 19180 36270 19220 36340
rect 19280 36270 19320 36340
rect 19380 36270 19420 36340
rect 19480 36270 19520 36340
rect 19580 36270 19620 36340
rect 19680 36270 19720 36340
rect 19780 36270 19820 36340
rect 19880 36270 19920 36340
rect 19980 36270 20020 36340
rect 20080 36270 20120 36340
rect 20180 36270 20220 36340
rect 20280 36270 20320 36340
rect 20380 36270 20420 36340
rect 20480 36270 20520 36340
rect 20580 36270 20620 36340
rect 20680 36270 20720 36340
rect 20780 36270 20820 36340
rect 20880 36270 20920 36340
rect 20980 36270 21020 36340
rect 21080 36270 21120 36340
rect 21180 36270 21220 36340
rect 21280 36270 21320 36340
rect 21380 36270 21420 36340
rect 21480 36270 21520 36340
rect 21580 36270 21620 36340
rect 21680 36270 21720 36340
rect 21780 36270 21820 36340
rect 21880 36270 21920 36340
rect 21980 36270 22020 36340
rect 22080 36270 22120 36340
rect 22180 36270 22220 36340
rect 22280 36270 22320 36340
rect 22380 36270 22420 36340
rect 22480 36270 22520 36340
rect 22580 36270 22620 36340
rect 22680 36270 22720 36340
rect 22780 36270 22820 36340
rect 22880 36270 22920 36340
rect 22980 36270 23020 36340
rect 23080 36270 23120 36340
rect 23180 36270 23220 36340
rect 23280 36270 23320 36340
rect 23380 36270 23420 36340
rect 23480 36270 23520 36340
rect 23580 36270 23620 36340
rect 23680 36270 23720 36340
rect 23780 36270 23820 36340
rect 23880 36270 23920 36340
rect 23980 36270 24020 36340
rect 24080 36270 24120 36340
rect 24180 36270 24220 36340
rect 24280 36270 24320 36340
rect 24380 36270 24420 36340
rect 24480 36270 24520 36340
rect 24580 36270 24620 36340
rect 24680 36270 24720 36340
rect 24780 36270 24820 36340
rect 24880 36270 24910 36340
rect 15180 36260 24910 36270
rect 15160 36110 15400 36120
rect 15160 36050 15200 36110
rect 15300 36050 15400 36110
rect 15440 36110 15520 36120
rect 15440 36070 15460 36110
rect 15500 36070 15520 36110
rect 15440 36060 15520 36070
rect 15160 36040 15400 36050
rect 15340 35950 15400 36040
rect 15340 35790 15350 35950
rect 15390 35790 15400 35950
rect 15340 35770 15400 35790
rect 15450 35950 15510 36060
rect 15450 35790 15460 35950
rect 15500 35790 15510 35950
rect 15450 35520 15510 35790
rect 15560 35950 15620 35970
rect 15560 35790 15570 35950
rect 15610 35790 15620 35950
rect 15560 35740 15620 35790
rect 16460 35820 16520 36260
rect 15560 35680 15870 35740
rect 15820 35640 15870 35680
rect 15550 35630 15660 35640
rect 15550 35570 15570 35630
rect 15640 35570 15660 35630
rect 15550 35560 15660 35570
rect 15760 35630 15930 35640
rect 15760 35570 15790 35630
rect 15900 35570 15930 35630
rect 16460 35630 16470 35820
rect 16510 35630 16520 35820
rect 16460 35610 16520 35630
rect 16570 35820 16630 35840
rect 16570 35630 16580 35820
rect 16620 35630 16630 35820
rect 15760 35560 15930 35570
rect 15450 35480 15460 35520
rect 15500 35480 15510 35520
rect 16570 35550 16630 35630
rect 16680 35820 16740 36260
rect 16680 35630 16690 35820
rect 16730 35630 16740 35820
rect 16680 35610 16740 35630
rect 16790 35820 16850 35840
rect 16790 35630 16800 35820
rect 16840 35630 16850 35820
rect 16790 35550 16850 35630
rect 16900 35820 16960 36260
rect 16900 35630 16910 35820
rect 16950 35630 16960 35820
rect 16900 35610 16960 35630
rect 17010 35820 17070 35840
rect 17010 35630 17020 35820
rect 17060 35630 17070 35820
rect 17010 35550 17070 35630
rect 17120 35820 17180 36260
rect 17120 35630 17130 35820
rect 17170 35630 17180 35820
rect 17120 35610 17180 35630
rect 17460 36060 17520 36080
rect 17460 35600 17470 36060
rect 17510 35600 17520 36060
rect 16570 35510 17200 35550
rect 15450 35460 15510 35480
rect 16430 35490 16530 35510
rect 16430 35430 16450 35490
rect 16510 35430 16530 35490
rect 17120 35490 17200 35510
rect 17120 35450 17140 35490
rect 17180 35450 17200 35490
rect 17120 35430 17200 35450
rect 16430 35410 16530 35430
rect 16570 35390 17200 35430
rect 16460 35330 16520 35350
rect 6450 34810 6640 34850
rect 6680 34810 6720 34850
rect 6760 34810 6770 34850
rect 6450 34800 6770 34810
rect 3770 34790 5300 34800
rect 3770 34670 3830 34790
rect 3770 33710 3780 34670
rect 3820 33710 3830 34670
rect 3770 33690 3830 33710
rect 3880 34670 3940 34690
rect 3880 33710 3890 34670
rect 3930 33710 3940 34670
rect 3880 33630 3940 33710
rect 3990 34670 4050 34790
rect 3990 33710 4000 34670
rect 4040 33710 4050 34670
rect 3990 33690 4050 33710
rect 4100 34670 4160 34690
rect 4100 33710 4110 34670
rect 4150 33710 4160 34670
rect 4100 33630 4160 33710
rect 4210 34670 4270 34790
rect 4210 33710 4220 34670
rect 4260 33710 4270 34670
rect 4210 33690 4270 33710
rect 4320 34670 4380 34690
rect 4320 33710 4330 34670
rect 4370 33710 4380 34670
rect 4320 33630 4380 33710
rect 4500 34670 4570 34790
rect 4500 33710 4510 34670
rect 4560 33710 4570 34670
rect 4500 33690 4570 33710
rect 4690 34670 4750 34690
rect 4690 33710 4700 34670
rect 4740 33710 4750 34670
rect 4690 33630 4750 33710
rect 4800 34670 4860 34790
rect 4800 33710 4810 34670
rect 4850 33710 4860 34670
rect 4800 33690 4860 33710
rect 4910 34670 4970 34690
rect 4910 33710 4920 34670
rect 4960 33710 4970 34670
rect 4910 33630 4970 33710
rect 5020 34670 5080 34790
rect 5020 33710 5030 34670
rect 5070 33710 5080 34670
rect 5020 33690 5080 33710
rect 5130 34670 5190 34690
rect 5130 33710 5140 34670
rect 5180 33710 5190 34670
rect 5130 33630 5190 33710
rect 5240 34670 5300 34790
rect 5240 33710 5250 34670
rect 5290 33710 5300 34670
rect 5460 34740 5520 34760
rect 5460 33780 5470 34740
rect 5510 33780 5520 34740
rect 5460 33760 5520 33780
rect 5570 34740 5630 34760
rect 5570 33780 5580 34740
rect 5620 33780 5630 34740
rect 5240 33690 5300 33710
rect 5570 33630 5630 33780
rect 5680 34740 5740 34760
rect 5680 33780 5690 34740
rect 5730 33780 5740 34740
rect 5680 33760 5740 33780
rect 5790 34740 5850 34760
rect 5790 33780 5800 34740
rect 5840 33780 5850 34740
rect 5790 33630 5850 33780
rect 5900 34740 5960 34760
rect 5900 33780 5910 34740
rect 5950 33780 5960 34740
rect 5900 33760 5960 33780
rect 6010 34740 6070 34760
rect 6010 33780 6020 34740
rect 6060 33780 6070 34740
rect 6010 33630 6070 33780
rect 6120 34740 6180 34800
rect 6120 33780 6130 34740
rect 6170 33780 6180 34740
rect 6340 34740 6400 34760
rect 6340 34280 6350 34740
rect 6390 34280 6400 34740
rect 6340 34050 6400 34280
rect 6450 34740 6510 34800
rect 6710 34790 6770 34800
rect 6940 34840 7370 34850
rect 6940 34800 7220 34840
rect 7260 34800 7300 34840
rect 7340 34800 7370 34840
rect 6940 34790 7370 34800
rect 7410 34840 7750 34850
rect 7410 34800 7600 34840
rect 7640 34800 7680 34840
rect 7720 34800 7750 34840
rect 7410 34790 7750 34800
rect 7790 34840 8130 34850
rect 7790 34800 7980 34840
rect 8020 34800 8060 34840
rect 8100 34800 8130 34840
rect 7790 34790 8130 34800
rect 8170 34840 8510 34850
rect 8170 34800 8360 34840
rect 8400 34800 8440 34840
rect 8480 34800 8510 34840
rect 8170 34790 8510 34800
rect 8550 34840 8850 34850
rect 8550 34800 8690 34840
rect 8730 34800 8800 34840
rect 8840 34800 8850 34840
rect 8550 34790 8850 34800
rect 6450 34280 6460 34740
rect 6500 34280 6510 34740
rect 6450 34260 6510 34280
rect 6560 34740 6620 34760
rect 6560 34280 6570 34740
rect 6610 34280 6620 34740
rect 6560 34050 6620 34280
rect 6810 34730 6870 34750
rect 6810 34270 6820 34730
rect 6860 34270 6870 34730
rect 6810 34050 6870 34270
rect 6940 34730 7000 34790
rect 6940 34270 6950 34730
rect 6990 34270 7000 34730
rect 6940 34250 7000 34270
rect 7070 34730 7130 34750
rect 7070 34270 7080 34730
rect 7120 34270 7130 34730
rect 7070 34050 7130 34270
rect 7300 34730 7360 34750
rect 7300 34270 7310 34730
rect 7350 34270 7360 34730
rect 7170 34190 7230 34210
rect 7170 34150 7180 34190
rect 7220 34150 7230 34190
rect 7170 34130 7230 34150
rect 7300 34050 7360 34270
rect 7410 34730 7470 34790
rect 7410 34270 7420 34730
rect 7460 34270 7470 34730
rect 7410 34250 7470 34270
rect 7520 34730 7580 34750
rect 7520 34270 7530 34730
rect 7570 34270 7580 34730
rect 7520 34050 7580 34270
rect 7680 34730 7740 34750
rect 7680 34270 7690 34730
rect 7730 34270 7740 34730
rect 7680 34050 7740 34270
rect 7790 34730 7850 34790
rect 7790 34270 7800 34730
rect 7840 34270 7850 34730
rect 7790 34250 7850 34270
rect 7900 34730 7960 34750
rect 7900 34270 7910 34730
rect 7950 34270 7960 34730
rect 7900 34050 7960 34270
rect 8060 34730 8120 34750
rect 8060 34270 8070 34730
rect 8110 34270 8120 34730
rect 8060 34050 8120 34270
rect 8170 34730 8230 34790
rect 8170 34270 8180 34730
rect 8220 34270 8230 34730
rect 8170 34250 8230 34270
rect 8280 34730 8340 34750
rect 8280 34270 8290 34730
rect 8330 34270 8340 34730
rect 8280 34050 8340 34270
rect 8440 34730 8500 34750
rect 8440 34270 8450 34730
rect 8490 34270 8500 34730
rect 8440 34050 8500 34270
rect 8550 34730 8610 34790
rect 8790 34780 8850 34790
rect 9020 34840 9450 34850
rect 9020 34800 9300 34840
rect 9340 34800 9380 34840
rect 9420 34800 9450 34840
rect 9020 34790 9450 34800
rect 9490 34840 9830 34850
rect 9490 34800 9680 34840
rect 9720 34800 9760 34840
rect 9800 34800 9830 34840
rect 9490 34790 9830 34800
rect 9870 34840 10210 34850
rect 9870 34800 10060 34840
rect 10100 34800 10140 34840
rect 10180 34800 10210 34840
rect 9870 34790 10210 34800
rect 10250 34840 10590 34850
rect 10250 34800 10440 34840
rect 10480 34800 10520 34840
rect 10560 34800 10590 34840
rect 10250 34790 10590 34800
rect 10630 34840 10880 34850
rect 10630 34800 10820 34840
rect 10860 34800 10880 34840
rect 10630 34790 10880 34800
rect 8550 34270 8560 34730
rect 8600 34270 8610 34730
rect 8550 34250 8610 34270
rect 8660 34730 8720 34750
rect 8660 34270 8670 34730
rect 8710 34270 8720 34730
rect 8660 34050 8720 34270
rect 8890 34730 8950 34750
rect 8890 34270 8900 34730
rect 8940 34270 8950 34730
rect 8890 34050 8950 34270
rect 9020 34730 9080 34790
rect 9020 34270 9030 34730
rect 9070 34270 9080 34730
rect 9020 34250 9080 34270
rect 9150 34730 9210 34750
rect 9150 34270 9160 34730
rect 9200 34270 9210 34730
rect 9150 34050 9210 34270
rect 9380 34730 9440 34750
rect 9380 34270 9390 34730
rect 9430 34270 9440 34730
rect 9380 34050 9440 34270
rect 9490 34730 9550 34790
rect 9490 34270 9500 34730
rect 9540 34270 9550 34730
rect 9490 34250 9550 34270
rect 9600 34730 9660 34750
rect 9600 34270 9610 34730
rect 9650 34270 9660 34730
rect 9600 34050 9660 34270
rect 9760 34730 9820 34750
rect 9760 34270 9770 34730
rect 9810 34270 9820 34730
rect 9760 34050 9820 34270
rect 9870 34730 9930 34790
rect 9870 34270 9880 34730
rect 9920 34270 9930 34730
rect 9870 34250 9930 34270
rect 9980 34730 10040 34750
rect 9980 34270 9990 34730
rect 10030 34270 10040 34730
rect 9980 34050 10040 34270
rect 10140 34730 10200 34750
rect 10140 34270 10150 34730
rect 10190 34270 10200 34730
rect 10140 34050 10200 34270
rect 10250 34730 10310 34790
rect 10250 34270 10260 34730
rect 10300 34270 10310 34730
rect 10250 34250 10310 34270
rect 10360 34730 10420 34750
rect 10360 34270 10370 34730
rect 10410 34270 10420 34730
rect 10360 34050 10420 34270
rect 10520 34730 10580 34750
rect 10520 34270 10530 34730
rect 10570 34270 10580 34730
rect 10520 34050 10580 34270
rect 10630 34730 10690 34790
rect 10630 34270 10640 34730
rect 10680 34270 10690 34730
rect 10630 34250 10690 34270
rect 10740 34730 10800 34750
rect 10740 34270 10750 34730
rect 10790 34270 10800 34730
rect 10740 34050 10800 34270
rect 16460 34470 16470 35330
rect 16510 34470 16520 35330
rect 16460 34210 16520 34470
rect 16570 35330 16630 35390
rect 16570 34470 16580 35330
rect 16620 34470 16630 35330
rect 16570 34450 16630 34470
rect 16680 35330 16740 35350
rect 16680 34470 16690 35330
rect 16730 34470 16740 35330
rect 16680 34210 16740 34470
rect 16790 35330 16850 35390
rect 16790 34470 16800 35330
rect 16840 34470 16850 35330
rect 16790 34450 16850 34470
rect 16900 35330 16960 35350
rect 16900 34470 16910 35330
rect 16950 34470 16960 35330
rect 16900 34210 16960 34470
rect 17010 35330 17070 35390
rect 17010 34470 17020 35330
rect 17060 34470 17070 35330
rect 17010 34450 17070 34470
rect 17120 35330 17180 35350
rect 17120 34470 17130 35330
rect 17170 34470 17180 35330
rect 17460 35340 17520 35600
rect 17570 36060 17630 36260
rect 17570 35600 17580 36060
rect 17620 35600 17630 36060
rect 17570 35580 17630 35600
rect 17710 36060 17770 36260
rect 17710 35600 17720 36060
rect 17760 35600 17770 36060
rect 17710 35580 17770 35600
rect 17820 36060 17880 36080
rect 17820 35600 17830 36060
rect 17870 35600 17880 36060
rect 17560 35490 17780 35500
rect 17560 35450 17580 35490
rect 17620 35450 17720 35490
rect 17760 35450 17780 35490
rect 17560 35440 17780 35450
rect 17820 35490 17880 35600
rect 18030 36060 18090 36260
rect 18030 35600 18040 36060
rect 18080 35600 18090 36060
rect 18030 35580 18090 35600
rect 18140 36060 18200 36080
rect 18140 35600 18150 36060
rect 18190 35600 18200 36060
rect 18020 35490 18100 35500
rect 17820 35450 18040 35490
rect 18080 35450 18100 35490
rect 17640 35360 17700 35440
rect 17640 35340 17650 35360
rect 17460 35320 17650 35340
rect 17690 35320 17700 35360
rect 17820 35320 17880 35450
rect 18020 35440 18100 35450
rect 17460 35300 17700 35320
rect 17350 35140 17410 35160
rect 17350 34980 17360 35140
rect 17400 34980 17410 35140
rect 17350 34770 17410 34980
rect 17460 35140 17520 35300
rect 17460 34980 17470 35140
rect 17510 34980 17520 35140
rect 17460 34960 17520 34980
rect 17750 35270 17880 35320
rect 18140 35270 18200 35600
rect 18400 36060 18460 36080
rect 18400 35600 18410 36060
rect 18450 35600 18460 36060
rect 18400 35340 18460 35600
rect 18510 36060 18570 36260
rect 18510 35600 18520 36060
rect 18560 35600 18570 36060
rect 18510 35580 18570 35600
rect 18650 36060 18710 36260
rect 18650 35600 18660 36060
rect 18700 35600 18710 36060
rect 18650 35580 18710 35600
rect 18760 36060 18820 36080
rect 18760 35600 18770 36060
rect 18810 35600 18820 36060
rect 18500 35490 18720 35500
rect 18500 35450 18520 35490
rect 18560 35450 18660 35490
rect 18700 35450 18720 35490
rect 18500 35440 18720 35450
rect 18760 35490 18820 35600
rect 18970 36060 19030 36260
rect 18970 35600 18980 36060
rect 19020 35600 19030 36060
rect 18970 35580 19030 35600
rect 19080 36060 19140 36080
rect 19080 35600 19090 36060
rect 19130 35600 19140 36060
rect 18960 35490 19040 35500
rect 18760 35450 18980 35490
rect 19020 35450 19040 35490
rect 18580 35360 18640 35440
rect 18580 35340 18590 35360
rect 18400 35320 18590 35340
rect 18630 35320 18640 35360
rect 18760 35320 18820 35450
rect 18960 35440 19040 35450
rect 18400 35300 18640 35320
rect 17750 35090 17810 35270
rect 18030 35210 18200 35270
rect 17850 35200 17930 35210
rect 17850 35160 17870 35200
rect 17910 35160 17930 35200
rect 17850 35150 17930 35160
rect 17750 34930 17760 35090
rect 17800 34930 17810 35090
rect 17750 34910 17810 34930
rect 17860 35090 17920 35110
rect 17860 34930 17870 35090
rect 17910 34930 17920 35090
rect 17450 34900 17530 34910
rect 17450 34860 17470 34900
rect 17510 34860 17530 34900
rect 17450 34850 17530 34860
rect 17860 34770 17920 34930
rect 17350 34710 17920 34770
rect 17120 34210 17180 34470
rect 17570 34620 17630 34640
rect 17570 34460 17580 34620
rect 17620 34460 17630 34620
rect 17570 34210 17630 34460
rect 17680 34620 17740 34710
rect 17680 34460 17690 34620
rect 17730 34460 17740 34620
rect 17680 34440 17740 34460
rect 18030 34620 18090 35210
rect 18290 35140 18350 35160
rect 18290 34980 18300 35140
rect 18340 34980 18350 35140
rect 18290 34770 18350 34980
rect 18400 35140 18460 35300
rect 18400 34980 18410 35140
rect 18450 34980 18460 35140
rect 18400 34960 18460 34980
rect 18690 35270 18820 35320
rect 19080 35270 19140 35600
rect 18690 35140 18750 35270
rect 18970 35210 19140 35270
rect 19300 35990 19360 36260
rect 19760 36080 19820 36260
rect 18690 34980 18700 35140
rect 18740 34980 18750 35140
rect 18690 34960 18750 34980
rect 18800 35140 18860 35160
rect 18800 34980 18810 35140
rect 18850 34980 18860 35140
rect 18390 34900 18470 34910
rect 18390 34860 18410 34900
rect 18450 34860 18470 34900
rect 18390 34850 18470 34860
rect 18680 34900 18760 34910
rect 18680 34860 18700 34900
rect 18740 34860 18760 34900
rect 18680 34850 18760 34860
rect 18800 34770 18860 34980
rect 18290 34710 18860 34770
rect 18970 34970 19030 35210
rect 19300 35030 19310 35990
rect 19350 35030 19360 35990
rect 19300 35010 19360 35030
rect 19410 35990 19470 36010
rect 19410 35030 19420 35990
rect 19460 35030 19470 35990
rect 19760 35620 19770 36080
rect 19810 35620 19820 36080
rect 19760 35600 19820 35620
rect 19870 36080 19930 36100
rect 19870 35620 19880 36080
rect 19920 35620 19930 36080
rect 19870 35530 19930 35620
rect 20010 36080 20070 36260
rect 20010 35620 20020 36080
rect 20060 35620 20070 36080
rect 20010 35600 20070 35620
rect 20120 36080 20180 36100
rect 20120 35620 20130 36080
rect 20170 35620 20180 36080
rect 21030 35990 21090 36260
rect 19870 35520 20080 35530
rect 19750 35490 19830 35500
rect 19750 35450 19770 35490
rect 19810 35450 19830 35490
rect 19750 35440 19830 35450
rect 19870 35480 20020 35520
rect 20060 35480 20080 35520
rect 19870 35470 20080 35480
rect 19410 34970 19470 35030
rect 19760 35130 19820 35150
rect 19760 34970 19770 35130
rect 19810 34970 19820 35130
rect 18970 34950 19200 34970
rect 18970 34910 19130 34950
rect 19170 34910 19200 34950
rect 18970 34890 19200 34910
rect 19310 34950 19370 34970
rect 19310 34910 19320 34950
rect 19360 34910 19370 34950
rect 19310 34890 19370 34910
rect 19410 34950 19580 34970
rect 19410 34910 19520 34950
rect 19560 34910 19580 34950
rect 19410 34890 19580 34910
rect 19760 34910 19820 34970
rect 19870 35130 19930 35470
rect 20120 35390 20180 35620
rect 20120 35370 20260 35390
rect 20120 35330 20210 35370
rect 20250 35330 20260 35370
rect 20120 35310 20260 35330
rect 19870 34970 19880 35130
rect 19920 34970 19930 35130
rect 19870 34950 19930 34970
rect 20010 35130 20070 35150
rect 20010 34970 20020 35130
rect 20060 34970 20070 35130
rect 20010 34910 20070 34970
rect 20120 35130 20180 35310
rect 20120 34970 20130 35130
rect 20170 34970 20180 35130
rect 21030 35030 21040 35990
rect 21080 35030 21090 35990
rect 21030 35010 21090 35030
rect 21140 35990 21200 36010
rect 21140 35030 21150 35990
rect 21190 35030 21200 35990
rect 21420 35820 21480 36260
rect 21420 35630 21430 35820
rect 21470 35630 21480 35820
rect 21420 35610 21480 35630
rect 21530 35820 21590 35840
rect 21530 35630 21540 35820
rect 21580 35630 21590 35820
rect 21530 35550 21590 35630
rect 21640 35820 21700 36260
rect 21640 35630 21650 35820
rect 21690 35630 21700 35820
rect 21640 35610 21700 35630
rect 21750 35820 21810 35840
rect 21750 35630 21760 35820
rect 21800 35630 21810 35820
rect 21750 35550 21810 35630
rect 21860 35820 21920 36260
rect 21860 35630 21870 35820
rect 21910 35630 21920 35820
rect 21860 35610 21920 35630
rect 21970 35820 22030 35840
rect 21970 35630 21980 35820
rect 22020 35630 22030 35820
rect 21970 35550 22030 35630
rect 22080 35820 22140 36260
rect 22080 35630 22090 35820
rect 22130 35630 22140 35820
rect 22080 35610 22140 35630
rect 22420 36060 22480 36080
rect 22420 35600 22430 36060
rect 22470 35600 22480 36060
rect 21530 35510 22160 35550
rect 21410 35490 21490 35500
rect 21410 35450 21430 35490
rect 21470 35450 21490 35490
rect 21410 35440 21490 35450
rect 22080 35490 22160 35510
rect 22080 35450 22100 35490
rect 22140 35450 22160 35490
rect 22080 35430 22160 35450
rect 21530 35390 22160 35430
rect 20120 34950 20180 34970
rect 20900 34960 21000 34980
rect 18030 34460 18040 34620
rect 18080 34460 18090 34620
rect 18030 34440 18090 34460
rect 18140 34620 18200 34640
rect 18510 34620 18570 34640
rect 18140 34460 18150 34620
rect 18190 34460 18200 34620
rect 17670 34360 18100 34370
rect 17670 34320 17690 34360
rect 17730 34320 17870 34360
rect 17910 34320 18040 34360
rect 18080 34320 18100 34360
rect 17670 34310 18100 34320
rect 18140 34210 18200 34460
rect 18510 34460 18520 34620
rect 18560 34460 18570 34620
rect 18510 34210 18570 34460
rect 18620 34620 18680 34710
rect 18620 34460 18630 34620
rect 18670 34460 18680 34620
rect 18620 34440 18680 34460
rect 18970 34620 19030 34890
rect 19300 34830 19360 34850
rect 18970 34460 18980 34620
rect 19020 34460 19030 34620
rect 18970 34440 19030 34460
rect 19080 34620 19140 34640
rect 19080 34460 19090 34620
rect 19130 34460 19140 34620
rect 18610 34360 19040 34370
rect 18610 34320 18630 34360
rect 18670 34320 18810 34360
rect 18850 34320 18980 34360
rect 19020 34320 19040 34360
rect 18610 34310 19040 34320
rect 19080 34210 19140 34460
rect 19300 34470 19310 34830
rect 19350 34470 19360 34830
rect 19300 34210 19360 34470
rect 19410 34830 19470 34890
rect 19760 34870 19930 34910
rect 19410 34470 19420 34830
rect 19460 34470 19470 34830
rect 19730 34810 19830 34830
rect 19730 34750 19750 34810
rect 19810 34750 19830 34810
rect 19730 34730 19830 34750
rect 19870 34820 19930 34870
rect 20010 34860 20180 34910
rect 20900 34900 20920 34960
rect 20980 34900 21000 34960
rect 20900 34880 21000 34900
rect 21140 34970 21200 35030
rect 21420 35330 21480 35350
rect 21140 34950 21240 34970
rect 21140 34910 21190 34950
rect 21230 34910 21240 34950
rect 21140 34890 21240 34910
rect 19870 34810 20080 34820
rect 19870 34770 19880 34810
rect 19920 34770 20020 34810
rect 20060 34770 20080 34810
rect 19870 34760 20080 34770
rect 19750 34660 19830 34670
rect 19750 34620 19770 34660
rect 19810 34620 19830 34660
rect 19750 34610 19830 34620
rect 19410 34450 19470 34470
rect 19760 34550 19820 34570
rect 19760 34390 19770 34550
rect 19810 34390 19820 34550
rect 19760 34210 19820 34390
rect 19870 34550 19930 34760
rect 19870 34390 19880 34550
rect 19920 34390 19930 34550
rect 19870 34370 19930 34390
rect 20120 34210 20180 34860
rect 21030 34830 21090 34850
rect 21030 34470 21040 34830
rect 21080 34470 21090 34830
rect 21030 34210 21090 34470
rect 21140 34830 21200 34890
rect 21140 34470 21150 34830
rect 21190 34470 21200 34830
rect 21140 34450 21200 34470
rect 21420 34470 21430 35330
rect 21470 34470 21480 35330
rect 21420 34210 21480 34470
rect 21530 35330 21590 35390
rect 21530 34470 21540 35330
rect 21580 34470 21590 35330
rect 21530 34450 21590 34470
rect 21640 35330 21700 35350
rect 21640 34470 21650 35330
rect 21690 34470 21700 35330
rect 21640 34210 21700 34470
rect 21750 35330 21810 35390
rect 21750 34470 21760 35330
rect 21800 34470 21810 35330
rect 21750 34450 21810 34470
rect 21860 35330 21920 35350
rect 21860 34470 21870 35330
rect 21910 34470 21920 35330
rect 21860 34210 21920 34470
rect 21970 35330 22030 35390
rect 21970 34470 21980 35330
rect 22020 34470 22030 35330
rect 21970 34450 22030 34470
rect 22080 35330 22140 35350
rect 22080 34470 22090 35330
rect 22130 34470 22140 35330
rect 22420 35340 22480 35600
rect 22530 36060 22590 36260
rect 22530 35600 22540 36060
rect 22580 35600 22590 36060
rect 22530 35580 22590 35600
rect 22670 36060 22730 36260
rect 22670 35600 22680 36060
rect 22720 35600 22730 36060
rect 22670 35580 22730 35600
rect 22780 36060 22840 36080
rect 22780 35600 22790 36060
rect 22830 35600 22840 36060
rect 22520 35490 22740 35500
rect 22520 35450 22540 35490
rect 22580 35450 22680 35490
rect 22720 35450 22740 35490
rect 22520 35440 22740 35450
rect 22780 35490 22840 35600
rect 22990 36060 23050 36260
rect 22990 35600 23000 36060
rect 23040 35600 23050 36060
rect 22990 35580 23050 35600
rect 23100 36060 23160 36080
rect 23100 35600 23110 36060
rect 23150 35600 23160 36060
rect 22980 35490 23060 35500
rect 22780 35450 23000 35490
rect 23040 35450 23060 35490
rect 22600 35360 22660 35440
rect 22600 35340 22610 35360
rect 22420 35320 22610 35340
rect 22650 35320 22660 35360
rect 22780 35320 22840 35450
rect 22980 35440 23060 35450
rect 22420 35300 22660 35320
rect 22310 35140 22370 35160
rect 22310 34980 22320 35140
rect 22360 34980 22370 35140
rect 22310 34770 22370 34980
rect 22420 35140 22480 35300
rect 22420 34980 22430 35140
rect 22470 34980 22480 35140
rect 22420 34960 22480 34980
rect 22710 35270 22840 35320
rect 23100 35270 23160 35600
rect 22710 35090 22770 35270
rect 22990 35210 23160 35270
rect 23360 36060 23420 36080
rect 23360 35600 23370 36060
rect 23410 35600 23420 36060
rect 23360 35340 23420 35600
rect 23470 36060 23530 36260
rect 23470 35600 23480 36060
rect 23520 35600 23530 36060
rect 23470 35580 23530 35600
rect 23610 36060 23670 36260
rect 23610 35600 23620 36060
rect 23660 35600 23670 36060
rect 23610 35580 23670 35600
rect 23720 36060 23780 36080
rect 23720 35600 23730 36060
rect 23770 35600 23780 36060
rect 23460 35490 23680 35500
rect 23460 35450 23480 35490
rect 23520 35450 23620 35490
rect 23660 35450 23680 35490
rect 23460 35440 23680 35450
rect 23720 35490 23780 35600
rect 23930 36060 23990 36260
rect 23930 35600 23940 36060
rect 23980 35600 23990 36060
rect 23930 35580 23990 35600
rect 24040 36060 24100 36080
rect 24040 35600 24050 36060
rect 24090 35600 24100 36060
rect 23920 35490 24000 35500
rect 23720 35450 23940 35490
rect 23980 35450 24000 35490
rect 23540 35360 23600 35440
rect 23540 35340 23550 35360
rect 23360 35320 23550 35340
rect 23590 35320 23600 35360
rect 23720 35320 23780 35450
rect 23920 35440 24000 35450
rect 23360 35300 23600 35320
rect 22810 35200 22890 35210
rect 22810 35160 22830 35200
rect 22870 35160 22890 35200
rect 22810 35150 22890 35160
rect 22710 34930 22720 35090
rect 22760 34930 22770 35090
rect 22710 34910 22770 34930
rect 22820 35090 22880 35110
rect 22820 34930 22830 35090
rect 22870 34930 22880 35090
rect 22410 34900 22490 34910
rect 22410 34860 22430 34900
rect 22470 34860 22490 34900
rect 22410 34850 22490 34860
rect 22820 34770 22880 34930
rect 22310 34710 22880 34770
rect 22080 34210 22140 34470
rect 22530 34620 22590 34640
rect 22530 34460 22540 34620
rect 22580 34460 22590 34620
rect 22530 34210 22590 34460
rect 22640 34620 22700 34710
rect 22640 34460 22650 34620
rect 22690 34460 22700 34620
rect 22640 34440 22700 34460
rect 22990 34620 23050 35210
rect 23250 35140 23310 35160
rect 23250 34980 23260 35140
rect 23300 34980 23310 35140
rect 23250 34770 23310 34980
rect 23360 35140 23420 35300
rect 23650 35270 23780 35320
rect 24040 35270 24100 35600
rect 23360 34980 23370 35140
rect 23410 34980 23420 35140
rect 23360 34960 23420 34980
rect 23650 35140 23710 35270
rect 23930 35210 24100 35270
rect 24260 35990 24320 36260
rect 24720 36080 24780 36260
rect 23650 34980 23660 35140
rect 23700 34980 23710 35140
rect 23650 34960 23710 34980
rect 23760 35140 23820 35160
rect 23760 34980 23770 35140
rect 23810 34980 23820 35140
rect 23350 34900 23430 34910
rect 23350 34860 23370 34900
rect 23410 34860 23430 34900
rect 23350 34850 23430 34860
rect 23640 34900 23720 34910
rect 23640 34860 23660 34900
rect 23700 34860 23720 34900
rect 23640 34850 23720 34860
rect 23760 34770 23820 34980
rect 23250 34710 23820 34770
rect 23930 34970 23990 35210
rect 24260 35030 24270 35990
rect 24310 35030 24320 35990
rect 24260 35010 24320 35030
rect 24370 35990 24430 36010
rect 24370 35030 24380 35990
rect 24420 35030 24430 35990
rect 24720 35620 24730 36080
rect 24770 35620 24780 36080
rect 24720 35600 24780 35620
rect 24830 36080 24890 36100
rect 24830 35620 24840 36080
rect 24880 35620 24890 36080
rect 24830 35530 24890 35620
rect 24970 36080 25030 36260
rect 24970 35620 24980 36080
rect 25020 35620 25030 36080
rect 24970 35600 25030 35620
rect 25080 36080 25140 36100
rect 25080 35620 25090 36080
rect 25130 35620 25140 36080
rect 24830 35520 25040 35530
rect 24710 35490 24790 35500
rect 24710 35450 24730 35490
rect 24770 35450 24790 35490
rect 24710 35440 24790 35450
rect 24830 35480 24980 35520
rect 25020 35480 25040 35520
rect 24830 35470 25040 35480
rect 24370 34970 24430 35030
rect 24720 35130 24780 35150
rect 24720 34970 24730 35130
rect 24770 34970 24780 35130
rect 23930 34950 24160 34970
rect 23930 34910 24090 34950
rect 24130 34910 24160 34950
rect 23930 34890 24160 34910
rect 24270 34950 24330 34970
rect 24270 34910 24280 34950
rect 24320 34910 24330 34950
rect 24270 34890 24330 34910
rect 24370 34950 24540 34970
rect 24370 34910 24480 34950
rect 24520 34910 24540 34950
rect 24370 34890 24540 34910
rect 24720 34910 24780 34970
rect 24830 35130 24890 35470
rect 25080 35390 25140 35620
rect 25080 35370 25220 35390
rect 25080 35330 25170 35370
rect 25210 35330 25220 35370
rect 25080 35310 25220 35330
rect 24830 34970 24840 35130
rect 24880 34970 24890 35130
rect 24830 34950 24890 34970
rect 24970 35130 25030 35150
rect 24970 34970 24980 35130
rect 25020 34970 25030 35130
rect 24970 34910 25030 34970
rect 25080 35130 25140 35310
rect 25080 34970 25090 35130
rect 25130 34970 25140 35130
rect 25080 34950 25140 34970
rect 22990 34460 23000 34620
rect 23040 34460 23050 34620
rect 22990 34440 23050 34460
rect 23100 34620 23160 34640
rect 23100 34460 23110 34620
rect 23150 34460 23160 34620
rect 23470 34620 23530 34640
rect 22630 34360 23060 34370
rect 22630 34320 22650 34360
rect 22690 34320 22830 34360
rect 22870 34320 23000 34360
rect 23040 34320 23060 34360
rect 22630 34310 23060 34320
rect 23100 34210 23160 34460
rect 23470 34460 23480 34620
rect 23520 34460 23530 34620
rect 23470 34210 23530 34460
rect 23580 34620 23640 34710
rect 23580 34460 23590 34620
rect 23630 34460 23640 34620
rect 23580 34440 23640 34460
rect 23930 34620 23990 34890
rect 24260 34830 24320 34850
rect 23930 34460 23940 34620
rect 23980 34460 23990 34620
rect 23930 34440 23990 34460
rect 24040 34620 24100 34640
rect 24040 34460 24050 34620
rect 24090 34460 24100 34620
rect 23570 34360 24000 34370
rect 23570 34320 23590 34360
rect 23630 34320 23770 34360
rect 23810 34320 23940 34360
rect 23980 34320 24000 34360
rect 23570 34310 24000 34320
rect 24040 34210 24100 34460
rect 24260 34470 24270 34830
rect 24310 34470 24320 34830
rect 24260 34210 24320 34470
rect 24370 34830 24430 34890
rect 24720 34870 24890 34910
rect 24370 34470 24380 34830
rect 24420 34470 24430 34830
rect 24690 34810 24790 34830
rect 24690 34750 24710 34810
rect 24770 34750 24790 34810
rect 24690 34730 24790 34750
rect 24830 34820 24890 34870
rect 24970 34860 25140 34910
rect 24830 34810 25040 34820
rect 24830 34770 24840 34810
rect 24880 34770 24980 34810
rect 25020 34770 25040 34810
rect 24830 34760 25040 34770
rect 24710 34660 24790 34670
rect 24710 34620 24730 34660
rect 24770 34620 24790 34660
rect 24710 34610 24790 34620
rect 24370 34450 24430 34470
rect 24720 34550 24780 34570
rect 24720 34390 24730 34550
rect 24770 34390 24780 34550
rect 24720 34210 24780 34390
rect 24830 34550 24890 34760
rect 24830 34390 24840 34550
rect 24880 34390 24890 34550
rect 24830 34370 24890 34390
rect 25080 34210 25140 34860
rect 16460 34200 25450 34210
rect 16460 34130 16510 34200
rect 16570 34130 16610 34200
rect 16670 34130 16710 34200
rect 16770 34130 16810 34200
rect 16870 34130 16910 34200
rect 16970 34130 17010 34200
rect 17070 34130 17110 34200
rect 17170 34130 17210 34200
rect 17270 34130 17310 34200
rect 17370 34130 17410 34200
rect 17470 34130 17510 34200
rect 17570 34130 17610 34200
rect 17670 34130 17710 34200
rect 17770 34130 17810 34200
rect 17870 34130 17910 34200
rect 17970 34130 18010 34200
rect 18070 34130 18110 34200
rect 18170 34130 18210 34200
rect 18270 34130 18310 34200
rect 18370 34130 18410 34200
rect 18470 34130 18510 34200
rect 18570 34130 18610 34200
rect 18670 34130 18710 34200
rect 18770 34130 18810 34200
rect 18870 34130 18910 34200
rect 18970 34130 19010 34200
rect 19070 34130 19110 34200
rect 19170 34130 19210 34200
rect 19270 34130 19310 34200
rect 19370 34130 19410 34200
rect 19470 34130 19510 34200
rect 19570 34130 19610 34200
rect 19670 34130 19710 34200
rect 19770 34130 19810 34200
rect 19870 34130 19910 34200
rect 19970 34130 20010 34200
rect 20070 34130 20110 34200
rect 20170 34130 20210 34200
rect 20270 34130 20310 34200
rect 20370 34130 20410 34200
rect 20470 34130 20510 34200
rect 20570 34130 20610 34200
rect 20670 34130 20710 34200
rect 20770 34130 20810 34200
rect 20870 34130 20910 34200
rect 20970 34130 21010 34200
rect 21070 34130 21110 34200
rect 21170 34130 21210 34200
rect 21270 34130 21310 34200
rect 21370 34130 21410 34200
rect 21470 34130 21510 34200
rect 21570 34130 21610 34200
rect 21670 34130 21710 34200
rect 21770 34130 21810 34200
rect 21870 34130 21910 34200
rect 21970 34130 22010 34200
rect 22070 34130 22110 34200
rect 22170 34130 22210 34200
rect 22270 34130 22310 34200
rect 22370 34130 22410 34200
rect 22470 34130 22510 34200
rect 22570 34130 22610 34200
rect 22670 34130 22710 34200
rect 22770 34130 22810 34200
rect 22870 34130 22910 34200
rect 22970 34130 23010 34200
rect 23070 34130 23110 34200
rect 23170 34130 23210 34200
rect 23270 34130 23310 34200
rect 23370 34130 23410 34200
rect 23470 34130 23510 34200
rect 23570 34130 23620 34200
rect 23680 34130 23720 34200
rect 23780 34130 23820 34200
rect 23880 34130 23920 34200
rect 23980 34130 24020 34200
rect 24080 34130 24120 34200
rect 24180 34130 24220 34200
rect 24280 34130 24320 34200
rect 24380 34130 24420 34200
rect 24480 34130 24520 34200
rect 24580 34130 24620 34200
rect 24680 34130 24720 34200
rect 24780 34130 24820 34200
rect 24880 34130 24920 34200
rect 24980 34130 25020 34200
rect 25080 34130 25120 34200
rect 25180 34130 25220 34200
rect 25280 34130 25320 34200
rect 25380 34130 25450 34200
rect 16460 34120 25450 34130
rect 6340 34040 10880 34050
rect 6340 33980 6380 34040
rect 6440 33980 6480 34040
rect 6540 33980 6580 34040
rect 6640 33980 6680 34040
rect 6740 33980 6780 34040
rect 6840 33980 6880 34040
rect 6940 33980 6980 34040
rect 7040 33980 7080 34040
rect 7140 33980 7180 34040
rect 7240 33980 7280 34040
rect 7340 33980 7380 34040
rect 7440 33980 7480 34040
rect 7540 33980 7580 34040
rect 7640 33980 7680 34040
rect 7740 33980 7780 34040
rect 7840 33980 7880 34040
rect 7940 33980 7980 34040
rect 8040 33980 8080 34040
rect 8140 33980 8180 34040
rect 8240 33980 8280 34040
rect 8340 33980 8380 34040
rect 8440 33980 8480 34040
rect 8540 33980 8580 34040
rect 8640 33980 8680 34040
rect 8740 33980 8780 34040
rect 8840 33980 8880 34040
rect 8940 33980 8980 34040
rect 9040 33980 9080 34040
rect 9140 33980 9180 34040
rect 9240 33980 9280 34040
rect 9340 33980 9380 34040
rect 9440 33980 9480 34040
rect 9540 33980 9580 34040
rect 9640 33980 9680 34040
rect 9740 33980 9780 34040
rect 9840 33980 9880 34040
rect 9940 33980 9980 34040
rect 10040 33980 10080 34040
rect 10140 33980 10180 34040
rect 10240 33980 10280 34040
rect 10340 33980 10380 34040
rect 10440 33980 10480 34040
rect 10540 33980 10580 34040
rect 10640 33980 10680 34040
rect 10740 33980 10780 34040
rect 10840 33980 10880 34040
rect 6340 33970 10880 33980
rect 6120 33760 6180 33780
rect 3770 33620 6210 33630
rect 3770 33560 3810 33620
rect 3870 33560 3910 33620
rect 3970 33560 4010 33620
rect 4070 33560 4110 33620
rect 4170 33560 4210 33620
rect 4270 33560 4310 33620
rect 4370 33560 4410 33620
rect 4470 33560 4510 33620
rect 4570 33560 4610 33620
rect 4670 33560 4710 33620
rect 4770 33560 4810 33620
rect 4870 33560 4910 33620
rect 4970 33560 5010 33620
rect 5070 33560 5110 33620
rect 5170 33560 5210 33620
rect 5270 33560 5310 33620
rect 5370 33560 5410 33620
rect 5470 33560 5510 33620
rect 5570 33560 5610 33620
rect 5670 33560 5710 33620
rect 5770 33560 5810 33620
rect 5870 33560 5910 33620
rect 5970 33560 6010 33620
rect 6070 33560 6110 33620
rect 6170 33560 6210 33620
rect 3770 33550 6210 33560
rect 13728 32460 13950 32480
rect 13728 32420 13768 32460
rect 13848 32420 13950 32460
rect 13728 32400 13950 32420
rect 13890 32310 13950 32400
rect 14098 32380 14178 32390
rect 14098 32340 14118 32380
rect 14158 32340 14178 32380
rect 14098 32330 14178 32340
rect 13888 32280 13950 32310
rect 13888 32220 13948 32280
rect 13888 32060 13898 32220
rect 13938 32060 13948 32220
rect 13888 32040 13948 32060
rect 13998 32220 14058 32240
rect 13998 32060 14008 32220
rect 14048 32060 14058 32220
rect 13998 31950 14058 32060
rect 14108 32220 14168 32330
rect 14108 32060 14118 32220
rect 14158 32060 14168 32220
rect 13988 31940 14068 31950
rect 13988 31900 14008 31940
rect 14048 31900 14068 31940
rect 13988 31890 14068 31900
rect 14108 31790 14168 32060
rect 14218 32220 14278 32240
rect 14218 32060 14228 32220
rect 14268 32060 14278 32220
rect 16030 32180 25410 32190
rect 16030 32110 16120 32180
rect 16180 32110 16220 32180
rect 16280 32110 16320 32180
rect 16380 32110 16420 32180
rect 16480 32110 16520 32180
rect 16580 32110 16620 32180
rect 16680 32110 16720 32180
rect 16780 32110 16820 32180
rect 16880 32110 16920 32180
rect 16980 32110 17020 32180
rect 17080 32110 17120 32180
rect 17180 32110 17220 32180
rect 17280 32110 17320 32180
rect 17380 32110 17420 32180
rect 17480 32110 17520 32180
rect 17580 32110 17620 32180
rect 17680 32110 17720 32180
rect 17780 32110 17820 32180
rect 17880 32110 17920 32180
rect 17980 32110 18020 32180
rect 18080 32110 18120 32180
rect 18180 32110 18220 32180
rect 18280 32110 18320 32180
rect 18380 32110 18420 32180
rect 18480 32110 18520 32180
rect 18580 32110 18620 32180
rect 18680 32110 18720 32180
rect 18780 32110 18820 32180
rect 18880 32110 18920 32180
rect 18980 32110 19020 32180
rect 19080 32110 19120 32180
rect 19180 32110 19220 32180
rect 19280 32110 19320 32180
rect 19380 32110 19420 32180
rect 19480 32110 19520 32180
rect 19580 32110 19620 32180
rect 19680 32110 19720 32180
rect 19780 32110 19820 32180
rect 19880 32110 19920 32180
rect 19980 32110 20020 32180
rect 20080 32110 20120 32180
rect 20180 32110 20220 32180
rect 20280 32110 20320 32180
rect 20380 32110 20420 32180
rect 20480 32110 20520 32180
rect 20580 32110 20620 32180
rect 20680 32110 20720 32180
rect 20780 32110 20820 32180
rect 20880 32110 20920 32180
rect 20980 32110 21020 32180
rect 21080 32110 21120 32180
rect 21180 32110 21220 32180
rect 21280 32110 21320 32180
rect 21380 32110 21420 32180
rect 21480 32110 21520 32180
rect 21580 32110 21620 32180
rect 21680 32110 21720 32180
rect 21780 32110 21820 32180
rect 21880 32110 21920 32180
rect 21980 32110 22020 32180
rect 22080 32110 22120 32180
rect 22180 32110 22220 32180
rect 22280 32110 22320 32180
rect 22380 32110 22420 32180
rect 22480 32110 22520 32180
rect 22580 32110 22620 32180
rect 22680 32110 22720 32180
rect 22780 32110 22820 32180
rect 22880 32110 22920 32180
rect 22980 32110 23020 32180
rect 23080 32110 23120 32180
rect 23180 32110 23220 32180
rect 23280 32110 23320 32180
rect 23380 32110 23420 32180
rect 23480 32110 23520 32180
rect 23580 32110 23620 32180
rect 23680 32110 23720 32180
rect 23780 32110 23820 32180
rect 23880 32110 23920 32180
rect 23980 32110 24020 32180
rect 24080 32110 24120 32180
rect 24180 32110 24220 32180
rect 24280 32110 24320 32180
rect 24380 32110 24420 32180
rect 24480 32110 24520 32180
rect 24580 32110 24620 32180
rect 24680 32110 24720 32180
rect 24780 32110 24820 32180
rect 24880 32110 24920 32180
rect 24980 32110 25020 32180
rect 25080 32110 25120 32180
rect 25180 32110 25220 32180
rect 25280 32110 25320 32180
rect 25380 32110 25410 32180
rect 16030 32100 25410 32110
rect 14218 32010 14278 32060
rect 14370 32010 14540 32020
rect 14218 31950 14400 32010
rect 14510 31950 14540 32010
rect 14370 31940 14540 31950
rect 14208 31890 14288 31900
rect 14208 31850 14228 31890
rect 14268 31850 14288 31890
rect 14208 31840 14288 31850
rect 14108 31750 14118 31790
rect 14158 31750 14168 31790
rect 14488 31780 14540 31940
rect 2170 31730 6310 31740
rect 2170 31670 2210 31730
rect 2270 31670 2310 31730
rect 2370 31670 2410 31730
rect 2470 31670 2510 31730
rect 2570 31670 2610 31730
rect 2670 31670 2710 31730
rect 2770 31670 2810 31730
rect 2870 31670 2910 31730
rect 2970 31670 3010 31730
rect 3070 31670 3110 31730
rect 3170 31670 3210 31730
rect 3270 31670 3310 31730
rect 3370 31670 3410 31730
rect 3470 31670 3510 31730
rect 3570 31670 3610 31730
rect 3670 31670 3710 31730
rect 3770 31670 3810 31730
rect 3870 31670 3910 31730
rect 3970 31670 4010 31730
rect 4070 31670 4110 31730
rect 4170 31670 4210 31730
rect 4270 31670 4310 31730
rect 4370 31670 4410 31730
rect 4470 31670 4510 31730
rect 4570 31670 4610 31730
rect 4670 31670 4710 31730
rect 4770 31670 4810 31730
rect 4870 31670 4910 31730
rect 4970 31670 5010 31730
rect 5070 31670 5110 31730
rect 5170 31670 5210 31730
rect 5270 31670 5310 31730
rect 5370 31670 5410 31730
rect 5470 31670 5510 31730
rect 5570 31670 5610 31730
rect 5670 31670 5710 31730
rect 5770 31670 5810 31730
rect 5870 31670 5910 31730
rect 5970 31670 6010 31730
rect 6070 31670 6110 31730
rect 6170 31670 6210 31730
rect 6270 31670 6310 31730
rect 2170 31660 6310 31670
rect 2170 31580 2230 31660
rect 2170 30820 2180 31580
rect 2220 30820 2230 31580
rect 2170 30800 2230 30820
rect 2280 31580 2340 31600
rect 2280 30820 2290 31580
rect 2330 30820 2340 31580
rect 2280 30800 2340 30820
rect 2390 31580 2450 31600
rect 2390 30820 2400 31580
rect 2440 30820 2450 31580
rect 2390 30800 2450 30820
rect 2500 31580 2560 31600
rect 2500 30820 2510 31580
rect 2550 30820 2560 31580
rect 2500 30800 2560 30820
rect 2610 31580 2670 31600
rect 2610 30820 2620 31580
rect 2660 30820 2670 31580
rect 2610 30800 2670 30820
rect 2720 31580 2780 31600
rect 2720 30820 2730 31580
rect 2770 30820 2780 31580
rect 2720 30800 2780 30820
rect 2900 31580 2960 31600
rect 2900 30820 2910 31580
rect 2950 30820 2960 31580
rect 2900 30800 2960 30820
rect 3090 31580 3150 31600
rect 3090 30820 3100 31580
rect 3140 30820 3150 31580
rect 3090 30800 3150 30820
rect 3200 31580 3260 31600
rect 3200 30820 3210 31580
rect 3250 30820 3260 31580
rect 3200 30800 3260 30820
rect 3310 31580 3370 31600
rect 3310 30820 3320 31580
rect 3360 30820 3370 31580
rect 3310 30800 3370 30820
rect 3420 31580 3480 31600
rect 3420 30820 3430 31580
rect 3470 30820 3480 31580
rect 3420 30800 3480 30820
rect 3530 31580 3590 31600
rect 3530 30820 3540 31580
rect 3580 30820 3590 31580
rect 3530 30800 3590 30820
rect 3640 31580 3700 31600
rect 3640 30820 3650 31580
rect 3690 30820 3700 31580
rect 3860 31580 3920 31600
rect 3860 31220 3870 31580
rect 3910 31220 3920 31580
rect 3860 31200 3920 31220
rect 3970 31580 4030 31660
rect 3970 31220 3980 31580
rect 4020 31220 4030 31580
rect 3970 31200 4030 31220
rect 4080 31580 4140 31600
rect 4080 31220 4090 31580
rect 4130 31220 4140 31580
rect 4080 31200 4140 31220
rect 4190 31580 4250 31660
rect 4190 31220 4200 31580
rect 4240 31220 4250 31580
rect 4190 31200 4250 31220
rect 4300 31580 4360 31600
rect 4300 31220 4310 31580
rect 4350 31220 4360 31580
rect 4300 31200 4360 31220
rect 4410 31580 4470 31660
rect 4410 31220 4420 31580
rect 4460 31220 4470 31580
rect 4410 31200 4470 31220
rect 4520 31580 4580 31600
rect 4520 31220 4530 31580
rect 4570 31220 4580 31580
rect 2130 30740 2240 30760
rect 2130 30690 2160 30740
rect 2210 30690 2240 30740
rect 2130 30670 2240 30690
rect 2930 30740 3050 30760
rect 2930 30680 2960 30740
rect 3020 30680 3050 30740
rect 2930 30670 3050 30680
rect 3640 30620 3700 30820
rect 4520 30620 4580 31220
rect 4720 31580 4780 31600
rect 4720 31220 4730 31580
rect 4770 31220 4780 31580
rect 4720 31200 4780 31220
rect 4830 31580 4890 31660
rect 4830 31220 4840 31580
rect 4880 31220 4890 31580
rect 4830 31200 4890 31220
rect 4940 31580 5000 31600
rect 4940 31220 4950 31580
rect 4990 31220 5000 31580
rect 4940 31200 5000 31220
rect 5050 31580 5110 31660
rect 5050 31220 5060 31580
rect 5100 31220 5110 31580
rect 5050 31200 5110 31220
rect 5160 31580 5220 31600
rect 5160 31220 5170 31580
rect 5210 31220 5220 31580
rect 5160 31200 5220 31220
rect 5270 31580 5330 31660
rect 5270 31220 5280 31580
rect 5320 31220 5330 31580
rect 5270 31200 5330 31220
rect 5380 31580 5440 31600
rect 5380 31220 5390 31580
rect 5430 31220 5440 31580
rect 5380 30620 5440 31220
rect 5580 31580 5640 31600
rect 5580 31220 5590 31580
rect 5630 31220 5640 31580
rect 5580 31200 5640 31220
rect 5690 31580 5750 31660
rect 5690 31220 5700 31580
rect 5740 31220 5750 31580
rect 5690 31200 5750 31220
rect 5800 31580 5860 31600
rect 5800 31220 5810 31580
rect 5850 31220 5860 31580
rect 5800 31200 5860 31220
rect 5910 31580 5970 31660
rect 5910 31220 5920 31580
rect 5960 31220 5970 31580
rect 5910 31200 5970 31220
rect 6020 31580 6080 31600
rect 6020 31220 6030 31580
rect 6070 31220 6080 31580
rect 6020 31200 6080 31220
rect 6130 31580 6190 31660
rect 14108 31640 14168 31750
rect 6130 31220 6140 31580
rect 6180 31220 6190 31580
rect 6130 31200 6190 31220
rect 6240 31580 6300 31600
rect 6240 31220 6250 31580
rect 6290 31220 6300 31580
rect 6380 31380 11240 31400
rect 6380 31320 6470 31380
rect 6530 31320 6580 31380
rect 6640 31320 6690 31380
rect 6750 31320 6800 31380
rect 6860 31320 6910 31380
rect 6970 31320 7020 31380
rect 7080 31320 7130 31380
rect 7190 31320 7240 31380
rect 7300 31320 7350 31380
rect 7410 31320 7460 31380
rect 7520 31320 7570 31380
rect 7630 31320 7680 31380
rect 7740 31320 7790 31380
rect 7850 31320 7900 31380
rect 7960 31320 8010 31380
rect 8070 31320 8120 31380
rect 8180 31320 8230 31380
rect 8290 31320 8340 31380
rect 8400 31320 8450 31380
rect 8510 31320 8560 31380
rect 8620 31320 8670 31380
rect 8730 31320 8780 31380
rect 8840 31320 8890 31380
rect 8950 31320 9000 31380
rect 9060 31320 9110 31380
rect 9170 31320 9220 31380
rect 9280 31320 9330 31380
rect 9390 31320 9440 31380
rect 9500 31320 9550 31380
rect 9610 31320 9660 31380
rect 9720 31320 9770 31380
rect 9830 31320 9880 31380
rect 9940 31320 9990 31380
rect 10050 31320 10100 31380
rect 10160 31320 10210 31380
rect 10270 31320 10320 31380
rect 10380 31320 10430 31380
rect 10490 31320 10540 31380
rect 10600 31320 10650 31380
rect 10710 31320 10760 31380
rect 10820 31320 10880 31380
rect 10940 31320 10990 31380
rect 11050 31320 11100 31380
rect 11160 31320 11240 31380
rect 14108 31380 14118 31640
rect 14158 31380 14168 31640
rect 14108 31360 14168 31380
rect 14218 31730 14540 31780
rect 16460 31760 16520 32100
rect 14218 31640 14278 31730
rect 14218 31380 14228 31640
rect 14268 31380 14278 31640
rect 16460 31570 16470 31760
rect 16510 31570 16520 31760
rect 16460 31550 16520 31570
rect 16570 31760 16630 31780
rect 16570 31570 16580 31760
rect 16620 31570 16630 31760
rect 16570 31490 16630 31570
rect 16680 31760 16740 32100
rect 16680 31570 16690 31760
rect 16730 31570 16740 31760
rect 16680 31550 16740 31570
rect 16790 31760 16850 31780
rect 16790 31570 16800 31760
rect 16840 31570 16850 31760
rect 16790 31490 16850 31570
rect 16900 31760 16960 32100
rect 16900 31570 16910 31760
rect 16950 31570 16960 31760
rect 16900 31550 16960 31570
rect 17010 31760 17070 31780
rect 17010 31570 17020 31760
rect 17060 31570 17070 31760
rect 17010 31490 17070 31570
rect 17120 31760 17180 32100
rect 17120 31570 17130 31760
rect 17170 31570 17180 31760
rect 17120 31550 17180 31570
rect 17460 32000 17520 32020
rect 17460 31540 17470 32000
rect 17510 31540 17520 32000
rect 14218 31360 14278 31380
rect 16430 31450 16530 31470
rect 16570 31450 17200 31490
rect 16430 31390 16450 31450
rect 16510 31390 16530 31450
rect 16430 31370 16530 31390
rect 17120 31430 17200 31450
rect 17120 31390 17140 31430
rect 17180 31390 17200 31430
rect 17120 31370 17200 31390
rect 16570 31330 17200 31370
rect 6380 31300 11240 31320
rect 6240 30720 6300 31220
rect 6400 31220 6460 31300
rect 6400 31060 6410 31220
rect 6450 31060 6460 31220
rect 6400 31040 6460 31060
rect 6510 31220 6570 31240
rect 6510 31060 6520 31220
rect 6560 31060 6570 31220
rect 6240 30710 6380 30720
rect 6510 30710 6570 31060
rect 6620 31220 6680 31300
rect 6620 31060 6630 31220
rect 6670 31060 6680 31220
rect 6620 31040 6680 31060
rect 6870 31220 6930 31300
rect 6870 30860 6880 31220
rect 6920 30860 6930 31220
rect 6870 30840 6930 30860
rect 7130 31220 7190 31240
rect 7130 30860 7140 31220
rect 7180 30860 7190 31220
rect 7360 31220 7420 31300
rect 7360 31060 7370 31220
rect 7410 31060 7420 31220
rect 7360 31040 7420 31060
rect 7470 31220 7530 31240
rect 7470 31060 7480 31220
rect 7520 31060 7530 31220
rect 6770 30710 6830 30720
rect 6240 30660 6310 30710
rect 6360 30700 6470 30710
rect 6360 30660 6400 30700
rect 6440 30660 6470 30700
rect 6240 30650 6470 30660
rect 6510 30700 6830 30710
rect 7130 30700 7190 30860
rect 7470 30700 7530 31060
rect 7580 31220 7640 31300
rect 7580 31060 7590 31220
rect 7630 31060 7640 31220
rect 7580 31040 7640 31060
rect 7740 31220 7800 31300
rect 7740 31060 7750 31220
rect 7790 31060 7800 31220
rect 7740 31040 7800 31060
rect 7850 31220 7910 31240
rect 7850 31060 7860 31220
rect 7900 31060 7910 31220
rect 7850 30700 7910 31060
rect 7960 31220 8020 31300
rect 7960 31060 7970 31220
rect 8010 31060 8020 31220
rect 7960 31040 8020 31060
rect 8120 31220 8180 31300
rect 8120 31060 8130 31220
rect 8170 31060 8180 31220
rect 8120 31040 8180 31060
rect 8230 31220 8290 31240
rect 8230 31060 8240 31220
rect 8280 31060 8290 31220
rect 8230 30700 8290 31060
rect 8340 31220 8400 31300
rect 8340 31060 8350 31220
rect 8390 31060 8400 31220
rect 8340 31040 8400 31060
rect 8500 31220 8560 31300
rect 8500 31060 8510 31220
rect 8550 31060 8560 31220
rect 8500 31040 8560 31060
rect 8610 31220 8670 31240
rect 8610 31060 8620 31220
rect 8660 31060 8670 31220
rect 8610 30700 8670 31060
rect 8720 31220 8780 31300
rect 8720 31060 8730 31220
rect 8770 31060 8780 31220
rect 8720 31040 8780 31060
rect 8950 31220 9010 31300
rect 8950 30860 8960 31220
rect 9000 30860 9010 31220
rect 8950 30840 9010 30860
rect 9210 31220 9270 31240
rect 9210 30860 9220 31220
rect 9260 30860 9270 31220
rect 9440 31220 9500 31300
rect 9440 31060 9450 31220
rect 9490 31060 9500 31220
rect 9440 31040 9500 31060
rect 9550 31220 9610 31240
rect 9550 31060 9560 31220
rect 9600 31060 9610 31220
rect 9110 30800 9170 30820
rect 9110 30760 9120 30800
rect 9160 30760 9170 30800
rect 9110 30740 9170 30760
rect 8850 30700 8910 30710
rect 9210 30700 9270 30860
rect 9550 30700 9610 31060
rect 9660 31220 9720 31300
rect 9660 31060 9670 31220
rect 9710 31060 9720 31220
rect 9660 31040 9720 31060
rect 9820 31220 9880 31300
rect 9820 31060 9830 31220
rect 9870 31060 9880 31220
rect 9820 31040 9880 31060
rect 9930 31220 9990 31240
rect 9930 31060 9940 31220
rect 9980 31060 9990 31220
rect 9930 30700 9990 31060
rect 10040 31220 10100 31300
rect 10040 31060 10050 31220
rect 10090 31060 10100 31220
rect 10040 31040 10100 31060
rect 10200 31220 10260 31300
rect 10200 31060 10210 31220
rect 10250 31060 10260 31220
rect 10200 31040 10260 31060
rect 10310 31220 10370 31240
rect 10310 31060 10320 31220
rect 10360 31060 10370 31220
rect 10310 30700 10370 31060
rect 10420 31220 10480 31300
rect 10420 31060 10430 31220
rect 10470 31060 10480 31220
rect 10420 31040 10480 31060
rect 10580 31220 10640 31300
rect 10580 31060 10590 31220
rect 10630 31060 10640 31220
rect 10580 31040 10640 31060
rect 10690 31220 10750 31240
rect 10690 31060 10700 31220
rect 10740 31060 10750 31220
rect 10690 30700 10750 31060
rect 10800 31220 10860 31300
rect 10800 31060 10810 31220
rect 10850 31060 10860 31220
rect 10800 31040 10860 31060
rect 10960 31220 11020 31300
rect 10960 31060 10970 31220
rect 11010 31060 11020 31220
rect 10960 31040 11020 31060
rect 11070 31220 11130 31240
rect 11070 31060 11080 31220
rect 11120 31060 11130 31220
rect 11070 30740 11130 31060
rect 11180 31220 11240 31300
rect 14098 31310 14178 31320
rect 14098 31270 14118 31310
rect 14158 31270 14178 31310
rect 14098 31260 14178 31270
rect 16460 31270 16520 31290
rect 11180 31060 11190 31220
rect 11230 31060 11240 31220
rect 11180 31040 11240 31060
rect 11070 30720 11320 30740
rect 6510 30660 6700 30700
rect 6740 30660 6780 30700
rect 6820 30660 6830 30700
rect 6510 30650 6830 30660
rect 2170 30610 3800 30620
rect 4520 30610 4790 30620
rect 2170 30600 3930 30610
rect 2170 30560 3730 30600
rect 3770 30560 3820 30600
rect 3860 30560 3930 30600
rect 2170 30550 3930 30560
rect 4520 30560 4590 30610
rect 4640 30560 4680 30610
rect 4730 30560 4790 30610
rect 4520 30550 4790 30560
rect 5380 30610 5650 30620
rect 5380 30560 5450 30610
rect 5500 30560 5540 30610
rect 5590 30560 5650 30610
rect 5380 30550 5650 30560
rect 2170 30540 3800 30550
rect 2170 30420 2230 30540
rect 2170 29460 2180 30420
rect 2220 29460 2230 30420
rect 2170 29440 2230 29460
rect 2280 30420 2340 30440
rect 2280 29460 2290 30420
rect 2330 29460 2340 30420
rect 2280 29380 2340 29460
rect 2390 30420 2450 30540
rect 2390 29460 2400 30420
rect 2440 29460 2450 30420
rect 2390 29440 2450 29460
rect 2500 30420 2560 30440
rect 2500 29460 2510 30420
rect 2550 29460 2560 30420
rect 2500 29380 2560 29460
rect 2610 30420 2670 30540
rect 2610 29460 2620 30420
rect 2660 29460 2670 30420
rect 2610 29440 2670 29460
rect 2720 30420 2780 30440
rect 2720 29460 2730 30420
rect 2770 29460 2780 30420
rect 2720 29380 2780 29460
rect 2900 30420 2970 30540
rect 2900 29460 2910 30420
rect 2960 29460 2970 30420
rect 2900 29440 2970 29460
rect 3090 30420 3150 30440
rect 3090 29460 3100 30420
rect 3140 29460 3150 30420
rect 3090 29380 3150 29460
rect 3200 30420 3260 30540
rect 3200 29460 3210 30420
rect 3250 29460 3260 30420
rect 3200 29440 3260 29460
rect 3310 30420 3370 30440
rect 3310 29460 3320 30420
rect 3360 29460 3370 30420
rect 3310 29380 3370 29460
rect 3420 30420 3480 30540
rect 3420 29460 3430 30420
rect 3470 29460 3480 30420
rect 3420 29440 3480 29460
rect 3530 30420 3590 30440
rect 3530 29460 3540 30420
rect 3580 29460 3590 30420
rect 3530 29380 3590 29460
rect 3640 30420 3700 30540
rect 3640 29460 3650 30420
rect 3690 29460 3700 30420
rect 3860 30490 3920 30510
rect 3860 29530 3870 30490
rect 3910 29530 3920 30490
rect 3860 29510 3920 29530
rect 3970 30490 4030 30510
rect 3970 29530 3980 30490
rect 4020 29530 4030 30490
rect 3640 29440 3700 29460
rect 3970 29380 4030 29530
rect 4080 30490 4140 30510
rect 4080 29530 4090 30490
rect 4130 29530 4140 30490
rect 4080 29510 4140 29530
rect 4190 30490 4250 30510
rect 4190 29530 4200 30490
rect 4240 29530 4250 30490
rect 4190 29380 4250 29530
rect 4300 30490 4360 30510
rect 4300 29530 4310 30490
rect 4350 29530 4360 30490
rect 4300 29510 4360 29530
rect 4410 30490 4470 30510
rect 4410 29530 4420 30490
rect 4460 29530 4470 30490
rect 4410 29380 4470 29530
rect 4520 30490 4580 30550
rect 4520 29530 4530 30490
rect 4570 29530 4580 30490
rect 4520 29510 4580 29530
rect 4720 30490 4780 30510
rect 4720 29530 4730 30490
rect 4770 29530 4780 30490
rect 4720 29510 4780 29530
rect 4830 30490 4890 30510
rect 4830 29530 4840 30490
rect 4880 29530 4890 30490
rect 4830 29380 4890 29530
rect 4940 30490 5000 30510
rect 4940 29530 4950 30490
rect 4990 29530 5000 30490
rect 4940 29510 5000 29530
rect 5050 30490 5110 30510
rect 5050 29530 5060 30490
rect 5100 29530 5110 30490
rect 5050 29380 5110 29530
rect 5160 30490 5220 30510
rect 5160 29530 5170 30490
rect 5210 29530 5220 30490
rect 5160 29510 5220 29530
rect 5270 30490 5330 30510
rect 5270 29530 5280 30490
rect 5320 29530 5330 30490
rect 5270 29380 5330 29530
rect 5380 30490 5440 30550
rect 5380 29530 5390 30490
rect 5430 29530 5440 30490
rect 5380 29510 5440 29530
rect 5580 30490 5640 30510
rect 5580 29530 5590 30490
rect 5630 29530 5640 30490
rect 5580 29510 5640 29530
rect 5690 30490 5750 30510
rect 5690 29530 5700 30490
rect 5740 29530 5750 30490
rect 5690 29380 5750 29530
rect 5800 30490 5860 30510
rect 5800 29530 5810 30490
rect 5850 29530 5860 30490
rect 5800 29510 5860 29530
rect 5910 30490 5970 30510
rect 5910 29530 5920 30490
rect 5960 29530 5970 30490
rect 5910 29380 5970 29530
rect 6020 30490 6080 30510
rect 6020 29530 6030 30490
rect 6070 29530 6080 30490
rect 6020 29510 6080 29530
rect 6130 30490 6190 30510
rect 6130 29530 6140 30490
rect 6180 29530 6190 30490
rect 6130 29380 6190 29530
rect 6240 30490 6300 30650
rect 6240 29530 6250 30490
rect 6290 29530 6300 30490
rect 6400 30590 6460 30610
rect 6400 30130 6410 30590
rect 6450 30130 6460 30590
rect 6400 29910 6460 30130
rect 6510 30590 6570 30650
rect 6770 30640 6830 30650
rect 7000 30690 7430 30700
rect 7000 30650 7280 30690
rect 7320 30650 7360 30690
rect 7400 30650 7430 30690
rect 7000 30640 7430 30650
rect 7470 30690 7810 30700
rect 7470 30650 7660 30690
rect 7700 30650 7740 30690
rect 7780 30650 7810 30690
rect 7470 30640 7810 30650
rect 7850 30690 8190 30700
rect 7850 30650 8040 30690
rect 8080 30650 8120 30690
rect 8160 30650 8190 30690
rect 7850 30640 8190 30650
rect 8230 30690 8570 30700
rect 8230 30650 8420 30690
rect 8460 30650 8500 30690
rect 8540 30650 8570 30690
rect 8230 30640 8570 30650
rect 8610 30690 8910 30700
rect 8610 30650 8750 30690
rect 8790 30650 8860 30690
rect 8900 30650 8910 30690
rect 8610 30640 8910 30650
rect 6510 30130 6520 30590
rect 6560 30130 6570 30590
rect 6510 30110 6570 30130
rect 6620 30590 6680 30610
rect 6620 30130 6630 30590
rect 6670 30130 6680 30590
rect 6620 29910 6680 30130
rect 6870 30580 6930 30600
rect 6870 30120 6880 30580
rect 6920 30120 6930 30580
rect 6870 29910 6930 30120
rect 7000 30580 7060 30640
rect 7000 30120 7010 30580
rect 7050 30120 7060 30580
rect 7000 30100 7060 30120
rect 7130 30580 7190 30600
rect 7130 30120 7140 30580
rect 7180 30120 7190 30580
rect 7130 29910 7190 30120
rect 7360 30580 7420 30600
rect 7360 30120 7370 30580
rect 7410 30120 7420 30580
rect 7230 30040 7290 30060
rect 7230 30000 7240 30040
rect 7280 30000 7290 30040
rect 7230 29980 7290 30000
rect 7360 29910 7420 30120
rect 7470 30580 7530 30640
rect 7470 30120 7480 30580
rect 7520 30120 7530 30580
rect 7470 30100 7530 30120
rect 7580 30580 7640 30600
rect 7580 30120 7590 30580
rect 7630 30120 7640 30580
rect 7580 29910 7640 30120
rect 7740 30580 7800 30600
rect 7740 30120 7750 30580
rect 7790 30120 7800 30580
rect 7740 29910 7800 30120
rect 7850 30580 7910 30640
rect 7850 30120 7860 30580
rect 7900 30120 7910 30580
rect 7850 30100 7910 30120
rect 7960 30580 8020 30600
rect 7960 30120 7970 30580
rect 8010 30120 8020 30580
rect 7960 29910 8020 30120
rect 8120 30580 8180 30600
rect 8120 30120 8130 30580
rect 8170 30120 8180 30580
rect 8120 29910 8180 30120
rect 8230 30580 8290 30640
rect 8230 30120 8240 30580
rect 8280 30120 8290 30580
rect 8230 30100 8290 30120
rect 8340 30580 8400 30600
rect 8340 30120 8350 30580
rect 8390 30120 8400 30580
rect 8340 29910 8400 30120
rect 8500 30580 8560 30600
rect 8500 30120 8510 30580
rect 8550 30120 8560 30580
rect 8500 29910 8560 30120
rect 8610 30580 8670 30640
rect 8850 30630 8910 30640
rect 9080 30690 9510 30700
rect 9080 30650 9360 30690
rect 9400 30650 9440 30690
rect 9480 30650 9510 30690
rect 9080 30640 9510 30650
rect 9550 30690 9890 30700
rect 9550 30650 9740 30690
rect 9780 30650 9820 30690
rect 9860 30650 9890 30690
rect 9550 30640 9890 30650
rect 9930 30690 10270 30700
rect 9930 30650 10120 30690
rect 10160 30650 10200 30690
rect 10240 30650 10270 30690
rect 9930 30640 10270 30650
rect 10310 30690 10650 30700
rect 10310 30650 10500 30690
rect 10540 30650 10580 30690
rect 10620 30650 10650 30690
rect 10310 30640 10650 30650
rect 10690 30690 11030 30700
rect 10690 30650 10880 30690
rect 10920 30650 10960 30690
rect 11000 30650 11030 30690
rect 10690 30640 11030 30650
rect 11070 30660 11240 30720
rect 11300 30660 11320 30720
rect 11070 30640 11320 30660
rect 8610 30120 8620 30580
rect 8660 30120 8670 30580
rect 8610 30100 8670 30120
rect 8720 30580 8780 30600
rect 8720 30120 8730 30580
rect 8770 30120 8780 30580
rect 8720 29910 8780 30120
rect 8950 30580 9010 30600
rect 8950 30120 8960 30580
rect 9000 30120 9010 30580
rect 8950 29910 9010 30120
rect 9080 30580 9140 30640
rect 9080 30120 9090 30580
rect 9130 30120 9140 30580
rect 9080 30100 9140 30120
rect 9210 30580 9270 30600
rect 9210 30120 9220 30580
rect 9260 30120 9270 30580
rect 9210 29910 9270 30120
rect 9440 30580 9500 30600
rect 9440 30120 9450 30580
rect 9490 30120 9500 30580
rect 9440 29910 9500 30120
rect 9550 30580 9610 30640
rect 9550 30120 9560 30580
rect 9600 30120 9610 30580
rect 9550 30100 9610 30120
rect 9660 30580 9720 30600
rect 9660 30120 9670 30580
rect 9710 30120 9720 30580
rect 9660 29910 9720 30120
rect 9820 30580 9880 30600
rect 9820 30120 9830 30580
rect 9870 30120 9880 30580
rect 9820 29910 9880 30120
rect 9930 30580 9990 30640
rect 9930 30120 9940 30580
rect 9980 30120 9990 30580
rect 9930 30100 9990 30120
rect 10040 30580 10100 30600
rect 10040 30120 10050 30580
rect 10090 30120 10100 30580
rect 10040 29910 10100 30120
rect 10200 30580 10260 30600
rect 10200 30120 10210 30580
rect 10250 30120 10260 30580
rect 10200 29910 10260 30120
rect 10310 30580 10370 30640
rect 10310 30120 10320 30580
rect 10360 30120 10370 30580
rect 10310 30100 10370 30120
rect 10420 30580 10480 30600
rect 10420 30120 10430 30580
rect 10470 30120 10480 30580
rect 10420 29910 10480 30120
rect 10580 30580 10640 30600
rect 10580 30120 10590 30580
rect 10630 30120 10640 30580
rect 10580 29910 10640 30120
rect 10690 30580 10750 30640
rect 10690 30120 10700 30580
rect 10740 30120 10750 30580
rect 10690 30100 10750 30120
rect 10800 30580 10860 30600
rect 10800 30120 10810 30580
rect 10850 30120 10860 30580
rect 10800 29910 10860 30120
rect 10960 30580 11020 30600
rect 10960 30120 10970 30580
rect 11010 30120 11020 30580
rect 10960 29910 11020 30120
rect 11070 30580 11130 30640
rect 11070 30120 11080 30580
rect 11120 30120 11130 30580
rect 11070 30100 11130 30120
rect 11180 30580 11240 30600
rect 11180 30120 11190 30580
rect 11230 30120 11240 30580
rect 16460 30410 16470 31270
rect 16510 30410 16520 31270
rect 16460 30140 16520 30410
rect 16570 31270 16630 31330
rect 16570 30410 16580 31270
rect 16620 30410 16630 31270
rect 16570 30390 16630 30410
rect 16680 31270 16740 31290
rect 16680 30410 16690 31270
rect 16730 30410 16740 31270
rect 16680 30140 16740 30410
rect 16790 31270 16850 31330
rect 16790 30410 16800 31270
rect 16840 30410 16850 31270
rect 16790 30390 16850 30410
rect 16900 31270 16960 31290
rect 16900 30410 16910 31270
rect 16950 30410 16960 31270
rect 16900 30140 16960 30410
rect 17010 31270 17070 31330
rect 17010 30410 17020 31270
rect 17060 30410 17070 31270
rect 17010 30390 17070 30410
rect 17120 31270 17180 31290
rect 17120 30410 17130 31270
rect 17170 30410 17180 31270
rect 17460 31280 17520 31540
rect 17570 32000 17630 32100
rect 17570 31540 17580 32000
rect 17620 31540 17630 32000
rect 17570 31520 17630 31540
rect 17710 32000 17770 32100
rect 17710 31540 17720 32000
rect 17760 31540 17770 32000
rect 17710 31520 17770 31540
rect 17820 32000 17880 32020
rect 17820 31540 17830 32000
rect 17870 31540 17880 32000
rect 17560 31430 17780 31440
rect 17560 31390 17580 31430
rect 17620 31390 17720 31430
rect 17760 31390 17780 31430
rect 17560 31380 17780 31390
rect 17820 31430 17880 31540
rect 18030 32000 18090 32100
rect 18030 31540 18040 32000
rect 18080 31540 18090 32000
rect 18030 31520 18090 31540
rect 18140 32000 18200 32020
rect 18140 31540 18150 32000
rect 18190 31540 18200 32000
rect 18020 31430 18100 31440
rect 17820 31390 18040 31430
rect 18080 31390 18100 31430
rect 17640 31300 17700 31380
rect 17640 31280 17650 31300
rect 17460 31260 17650 31280
rect 17690 31260 17700 31300
rect 17820 31260 17880 31390
rect 18020 31380 18100 31390
rect 17460 31240 17700 31260
rect 17350 31080 17410 31100
rect 17350 30920 17360 31080
rect 17400 30920 17410 31080
rect 17350 30710 17410 30920
rect 17460 31080 17520 31240
rect 17460 30920 17470 31080
rect 17510 30920 17520 31080
rect 17460 30900 17520 30920
rect 17750 31210 17880 31260
rect 18140 31210 18200 31540
rect 17750 31030 17810 31210
rect 18030 31150 18200 31210
rect 18400 32000 18460 32020
rect 18400 31540 18410 32000
rect 18450 31540 18460 32000
rect 18400 31280 18460 31540
rect 18510 32000 18570 32100
rect 18510 31540 18520 32000
rect 18560 31540 18570 32000
rect 18510 31520 18570 31540
rect 18650 32000 18710 32100
rect 18650 31540 18660 32000
rect 18700 31540 18710 32000
rect 18650 31520 18710 31540
rect 18760 32000 18820 32020
rect 18760 31540 18770 32000
rect 18810 31540 18820 32000
rect 18500 31430 18720 31440
rect 18500 31390 18520 31430
rect 18560 31390 18660 31430
rect 18700 31390 18720 31430
rect 18500 31380 18720 31390
rect 18760 31430 18820 31540
rect 18970 32000 19030 32100
rect 18970 31540 18980 32000
rect 19020 31540 19030 32000
rect 18970 31520 19030 31540
rect 19080 32000 19140 32020
rect 19080 31540 19090 32000
rect 19130 31540 19140 32000
rect 18960 31430 19040 31440
rect 18760 31390 18980 31430
rect 19020 31390 19040 31430
rect 18580 31300 18640 31380
rect 18580 31280 18590 31300
rect 18400 31260 18590 31280
rect 18630 31260 18640 31300
rect 18760 31260 18820 31390
rect 18960 31380 19040 31390
rect 18400 31240 18640 31260
rect 17850 31140 17930 31150
rect 17850 31100 17870 31140
rect 17910 31100 17930 31140
rect 17850 31090 17930 31100
rect 17750 30870 17760 31030
rect 17800 30870 17810 31030
rect 17750 30850 17810 30870
rect 17860 31030 17920 31050
rect 17860 30870 17870 31030
rect 17910 30870 17920 31030
rect 17450 30840 17530 30850
rect 17450 30800 17470 30840
rect 17510 30800 17530 30840
rect 17450 30790 17530 30800
rect 17860 30710 17920 30870
rect 17350 30650 17920 30710
rect 17120 30140 17180 30410
rect 17570 30560 17630 30580
rect 17570 30400 17580 30560
rect 17620 30400 17630 30560
rect 17570 30140 17630 30400
rect 17680 30560 17740 30650
rect 17680 30400 17690 30560
rect 17730 30400 17740 30560
rect 17680 30380 17740 30400
rect 18030 30560 18090 31150
rect 18290 31080 18350 31100
rect 18290 30920 18300 31080
rect 18340 30920 18350 31080
rect 18290 30710 18350 30920
rect 18400 31080 18460 31240
rect 18690 31210 18820 31260
rect 19080 31210 19140 31540
rect 18690 31080 18750 31210
rect 18970 31150 19140 31210
rect 19300 31930 19360 32100
rect 18400 30920 18410 31080
rect 18450 30920 18460 31080
rect 18400 30900 18460 30920
rect 18690 30920 18700 31080
rect 18740 30920 18750 31080
rect 18690 30900 18750 30920
rect 18800 31080 18860 31100
rect 18800 30920 18810 31080
rect 18850 30920 18860 31080
rect 18390 30840 18470 30850
rect 18390 30800 18410 30840
rect 18450 30800 18470 30840
rect 18390 30790 18470 30800
rect 18680 30840 18760 30850
rect 18680 30800 18700 30840
rect 18740 30800 18760 30840
rect 18680 30790 18760 30800
rect 18800 30710 18860 30920
rect 18290 30650 18860 30710
rect 18970 30910 19030 31150
rect 19300 30970 19310 31930
rect 19350 30970 19360 31930
rect 19300 30950 19360 30970
rect 19410 31930 19470 31950
rect 19410 30970 19420 31930
rect 19460 30970 19470 31930
rect 19410 30910 19470 30970
rect 19560 31930 19620 32100
rect 20020 32000 20080 32100
rect 19560 30970 19570 31930
rect 19610 30970 19620 31930
rect 19560 30950 19620 30970
rect 19670 31930 19730 31950
rect 19670 30970 19680 31930
rect 19720 30970 19730 31930
rect 20020 31540 20030 32000
rect 20070 31540 20080 32000
rect 20020 31520 20080 31540
rect 20130 32000 20190 32020
rect 20130 31540 20140 32000
rect 20180 31540 20190 32000
rect 20130 31450 20190 31540
rect 20270 32000 20330 32100
rect 20270 31540 20280 32000
rect 20320 31540 20330 32000
rect 20270 31520 20330 31540
rect 20380 32000 20440 32020
rect 20380 31540 20390 32000
rect 20430 31540 20440 32000
rect 20130 31440 20340 31450
rect 20010 31430 20090 31440
rect 20010 31390 20030 31430
rect 20070 31390 20090 31430
rect 20010 31380 20090 31390
rect 20130 31400 20280 31440
rect 20320 31400 20340 31440
rect 20130 31390 20340 31400
rect 19670 30910 19730 30970
rect 20020 31070 20080 31090
rect 20020 30910 20030 31070
rect 20070 30910 20080 31070
rect 18970 30890 19200 30910
rect 18970 30850 19130 30890
rect 19170 30850 19200 30890
rect 18970 30830 19200 30850
rect 19310 30890 19370 30910
rect 19310 30850 19320 30890
rect 19360 30850 19370 30890
rect 19310 30830 19370 30850
rect 19410 30890 19520 30910
rect 19410 30850 19460 30890
rect 19500 30850 19520 30890
rect 19410 30830 19520 30850
rect 19570 30890 19630 30910
rect 19570 30850 19580 30890
rect 19620 30850 19630 30890
rect 19570 30830 19630 30850
rect 19670 30890 19840 30910
rect 19670 30850 19780 30890
rect 19820 30850 19840 30890
rect 19670 30830 19840 30850
rect 20020 30850 20080 30910
rect 20130 31070 20190 31390
rect 20380 31260 20440 31540
rect 21090 31930 21150 32100
rect 20380 31240 20520 31260
rect 20380 31200 20470 31240
rect 20510 31200 20520 31240
rect 20380 31180 20520 31200
rect 20130 30910 20140 31070
rect 20180 30910 20190 31070
rect 20130 30890 20190 30910
rect 20270 31070 20330 31090
rect 20270 30910 20280 31070
rect 20320 30910 20330 31070
rect 20270 30850 20330 30910
rect 20380 31070 20440 31180
rect 20380 30910 20390 31070
rect 20430 30910 20440 31070
rect 21090 30970 21100 31930
rect 21140 30970 21150 31930
rect 21090 30950 21150 30970
rect 21200 31930 21260 31950
rect 21200 30970 21210 31930
rect 21250 30970 21260 31930
rect 21480 31750 21540 32100
rect 21480 31560 21490 31750
rect 21530 31560 21540 31750
rect 21480 31540 21540 31560
rect 21590 31750 21650 31770
rect 21590 31560 21600 31750
rect 21640 31560 21650 31750
rect 21590 31480 21650 31560
rect 21700 31750 21760 32100
rect 21700 31560 21710 31750
rect 21750 31560 21760 31750
rect 21700 31540 21760 31560
rect 21810 31750 21870 31770
rect 21810 31560 21820 31750
rect 21860 31560 21870 31750
rect 21810 31480 21870 31560
rect 21920 31750 21980 32100
rect 21920 31560 21930 31750
rect 21970 31560 21980 31750
rect 21920 31540 21980 31560
rect 22030 31750 22090 31770
rect 22030 31560 22040 31750
rect 22080 31560 22090 31750
rect 22030 31480 22090 31560
rect 22140 31750 22200 32100
rect 22140 31560 22150 31750
rect 22190 31560 22200 31750
rect 22140 31540 22200 31560
rect 22480 31990 22540 32010
rect 22480 31530 22490 31990
rect 22530 31530 22540 31990
rect 21590 31440 22220 31480
rect 21470 31420 21550 31430
rect 21470 31380 21490 31420
rect 21530 31380 21550 31420
rect 21470 31370 21550 31380
rect 22140 31420 22220 31440
rect 22140 31380 22160 31420
rect 22200 31380 22220 31420
rect 22140 31360 22220 31380
rect 21590 31320 22220 31360
rect 20380 30890 20440 30910
rect 20960 30900 21060 30920
rect 18030 30400 18040 30560
rect 18080 30400 18090 30560
rect 18030 30380 18090 30400
rect 18140 30560 18200 30580
rect 18140 30400 18150 30560
rect 18190 30400 18200 30560
rect 18510 30560 18570 30580
rect 18510 30400 18520 30560
rect 18560 30400 18570 30560
rect 17670 30300 18100 30310
rect 17670 30260 17690 30300
rect 17730 30260 17870 30300
rect 17910 30260 18040 30300
rect 18080 30260 18100 30300
rect 17670 30250 18100 30260
rect 18140 30140 18200 30400
rect 18510 30140 18570 30400
rect 18620 30560 18680 30650
rect 18620 30400 18630 30560
rect 18670 30400 18680 30560
rect 18620 30380 18680 30400
rect 18970 30560 19030 30830
rect 19300 30770 19360 30790
rect 18970 30400 18980 30560
rect 19020 30400 19030 30560
rect 18970 30380 19030 30400
rect 19080 30560 19140 30580
rect 19080 30400 19090 30560
rect 19130 30400 19140 30560
rect 18610 30300 19040 30310
rect 18610 30260 18630 30300
rect 18670 30260 18810 30300
rect 18850 30260 18980 30300
rect 19020 30260 19040 30300
rect 18610 30250 19040 30260
rect 19080 30140 19140 30400
rect 19300 30410 19310 30770
rect 19350 30410 19360 30770
rect 19300 30140 19360 30410
rect 19410 30770 19470 30830
rect 19410 30410 19420 30770
rect 19460 30410 19470 30770
rect 19410 30390 19470 30410
rect 19560 30770 19620 30790
rect 19560 30410 19570 30770
rect 19610 30410 19620 30770
rect 19560 30140 19620 30410
rect 19670 30770 19730 30830
rect 20020 30810 20190 30850
rect 19670 30410 19680 30770
rect 19720 30410 19730 30770
rect 19990 30750 20090 30770
rect 19990 30690 20010 30750
rect 20070 30690 20090 30750
rect 19990 30670 20090 30690
rect 20130 30760 20190 30810
rect 20270 30800 20440 30850
rect 20960 30840 20980 30900
rect 21040 30840 21060 30900
rect 20130 30750 20340 30760
rect 20130 30710 20140 30750
rect 20180 30710 20280 30750
rect 20320 30710 20340 30750
rect 20130 30700 20340 30710
rect 20010 30600 20090 30610
rect 20010 30560 20030 30600
rect 20070 30560 20090 30600
rect 20010 30550 20090 30560
rect 19670 30390 19730 30410
rect 20020 30490 20080 30510
rect 20020 30330 20030 30490
rect 20070 30330 20080 30490
rect 20020 30140 20080 30330
rect 20130 30490 20190 30700
rect 20130 30330 20140 30490
rect 20180 30330 20190 30490
rect 20130 30310 20190 30330
rect 20380 30140 20440 30800
rect 20960 30820 21060 30840
rect 21200 30910 21260 30970
rect 21480 31260 21540 31280
rect 21200 30890 21300 30910
rect 21200 30850 21250 30890
rect 21290 30850 21300 30890
rect 21200 30830 21300 30850
rect 21090 30770 21150 30790
rect 21090 30410 21100 30770
rect 21140 30410 21150 30770
rect 21090 30140 21150 30410
rect 21200 30770 21260 30830
rect 21200 30410 21210 30770
rect 21250 30410 21260 30770
rect 21200 30390 21260 30410
rect 21480 30400 21490 31260
rect 21530 30400 21540 31260
rect 21480 30140 21540 30400
rect 21590 31260 21650 31320
rect 21590 30400 21600 31260
rect 21640 30400 21650 31260
rect 21590 30380 21650 30400
rect 21700 31260 21760 31280
rect 21700 30400 21710 31260
rect 21750 30400 21760 31260
rect 21700 30140 21760 30400
rect 21810 31260 21870 31320
rect 21810 30400 21820 31260
rect 21860 30400 21870 31260
rect 21810 30380 21870 30400
rect 21920 31260 21980 31280
rect 21920 30400 21930 31260
rect 21970 30400 21980 31260
rect 21920 30140 21980 30400
rect 22030 31260 22090 31320
rect 22030 30400 22040 31260
rect 22080 30400 22090 31260
rect 22030 30380 22090 30400
rect 22140 31260 22200 31280
rect 22140 30400 22150 31260
rect 22190 30400 22200 31260
rect 22480 31270 22540 31530
rect 22590 31990 22650 32100
rect 22590 31530 22600 31990
rect 22640 31530 22650 31990
rect 22590 31510 22650 31530
rect 22730 31990 22790 32100
rect 22730 31530 22740 31990
rect 22780 31530 22790 31990
rect 22730 31510 22790 31530
rect 22840 31990 22900 32010
rect 22840 31530 22850 31990
rect 22890 31530 22900 31990
rect 22580 31420 22800 31430
rect 22580 31380 22600 31420
rect 22640 31380 22740 31420
rect 22780 31380 22800 31420
rect 22580 31370 22800 31380
rect 22840 31420 22900 31530
rect 23050 31990 23110 32100
rect 23050 31530 23060 31990
rect 23100 31530 23110 31990
rect 23050 31510 23110 31530
rect 23160 31990 23220 32010
rect 23160 31530 23170 31990
rect 23210 31530 23220 31990
rect 23040 31420 23120 31430
rect 22840 31380 23060 31420
rect 23100 31380 23120 31420
rect 22660 31290 22720 31370
rect 22660 31270 22670 31290
rect 22480 31250 22670 31270
rect 22710 31250 22720 31290
rect 22840 31250 22900 31380
rect 23040 31370 23120 31380
rect 22480 31230 22720 31250
rect 22370 31070 22430 31090
rect 22370 30910 22380 31070
rect 22420 30910 22430 31070
rect 22370 30700 22430 30910
rect 22480 31070 22540 31230
rect 22480 30910 22490 31070
rect 22530 30910 22540 31070
rect 22480 30890 22540 30910
rect 22770 31200 22900 31250
rect 23160 31200 23220 31530
rect 22770 31020 22830 31200
rect 23050 31140 23220 31200
rect 23420 31990 23480 32010
rect 23420 31530 23430 31990
rect 23470 31530 23480 31990
rect 23420 31270 23480 31530
rect 23530 31990 23590 32100
rect 23530 31530 23540 31990
rect 23580 31530 23590 31990
rect 23530 31510 23590 31530
rect 23670 31990 23730 32100
rect 23670 31530 23680 31990
rect 23720 31530 23730 31990
rect 23670 31510 23730 31530
rect 23780 31990 23840 32010
rect 23780 31530 23790 31990
rect 23830 31530 23840 31990
rect 23520 31420 23740 31430
rect 23520 31380 23540 31420
rect 23580 31380 23680 31420
rect 23720 31380 23740 31420
rect 23520 31370 23740 31380
rect 23780 31420 23840 31530
rect 23990 31990 24050 32100
rect 23990 31530 24000 31990
rect 24040 31530 24050 31990
rect 23990 31510 24050 31530
rect 24100 31990 24160 32010
rect 24100 31530 24110 31990
rect 24150 31530 24160 31990
rect 23980 31420 24060 31430
rect 23780 31380 24000 31420
rect 24040 31380 24060 31420
rect 23600 31290 23660 31370
rect 23600 31270 23610 31290
rect 23420 31250 23610 31270
rect 23650 31250 23660 31290
rect 23780 31250 23840 31380
rect 23980 31370 24060 31380
rect 23420 31230 23660 31250
rect 22870 31130 22950 31140
rect 22870 31090 22890 31130
rect 22930 31090 22950 31130
rect 22870 31080 22950 31090
rect 22770 30860 22780 31020
rect 22820 30860 22830 31020
rect 22770 30840 22830 30860
rect 22880 31020 22940 31040
rect 22880 30860 22890 31020
rect 22930 30860 22940 31020
rect 22470 30830 22550 30840
rect 22470 30790 22490 30830
rect 22530 30790 22550 30830
rect 22470 30780 22550 30790
rect 22880 30700 22940 30860
rect 22370 30640 22940 30700
rect 22140 30140 22200 30400
rect 22590 30550 22650 30570
rect 22590 30390 22600 30550
rect 22640 30390 22650 30550
rect 22590 30140 22650 30390
rect 22700 30550 22760 30640
rect 22700 30390 22710 30550
rect 22750 30390 22760 30550
rect 22700 30370 22760 30390
rect 23050 30550 23110 31140
rect 23310 31070 23370 31090
rect 23310 30910 23320 31070
rect 23360 30910 23370 31070
rect 23310 30700 23370 30910
rect 23420 31070 23480 31230
rect 23710 31200 23840 31250
rect 24100 31200 24160 31530
rect 23420 30910 23430 31070
rect 23470 30910 23480 31070
rect 23420 30890 23480 30910
rect 23710 31070 23770 31200
rect 23990 31140 24160 31200
rect 24320 31920 24380 32100
rect 23710 30910 23720 31070
rect 23760 30910 23770 31070
rect 23710 30890 23770 30910
rect 23820 31070 23880 31090
rect 23820 30910 23830 31070
rect 23870 30910 23880 31070
rect 23410 30830 23490 30840
rect 23410 30790 23430 30830
rect 23470 30790 23490 30830
rect 23410 30780 23490 30790
rect 23700 30830 23780 30840
rect 23700 30790 23720 30830
rect 23760 30790 23780 30830
rect 23700 30780 23780 30790
rect 23820 30700 23880 30910
rect 23310 30640 23880 30700
rect 23990 30900 24050 31140
rect 24320 30960 24330 31920
rect 24370 30960 24380 31920
rect 24320 30940 24380 30960
rect 24430 31920 24490 31940
rect 24430 30960 24440 31920
rect 24480 30960 24490 31920
rect 24430 30900 24490 30960
rect 24580 31920 24640 32100
rect 24980 32010 25040 32100
rect 24580 30960 24590 31920
rect 24630 30960 24640 31920
rect 24580 30940 24640 30960
rect 24690 31920 24750 31940
rect 24690 30960 24700 31920
rect 24740 30960 24750 31920
rect 24980 31550 24990 32010
rect 25030 31550 25040 32010
rect 24980 31530 25040 31550
rect 25090 32010 25150 32030
rect 25090 31550 25100 32010
rect 25140 31550 25150 32010
rect 25090 31460 25150 31550
rect 25230 32010 25290 32100
rect 25230 31550 25240 32010
rect 25280 31550 25290 32010
rect 25230 31530 25290 31550
rect 25340 32010 25400 32030
rect 25340 31550 25350 32010
rect 25390 31550 25400 32010
rect 25090 31450 25300 31460
rect 24970 31420 25050 31430
rect 24970 31380 24990 31420
rect 25030 31380 25050 31420
rect 24970 31370 25050 31380
rect 25090 31410 25240 31450
rect 25280 31410 25300 31450
rect 25090 31400 25300 31410
rect 24690 30900 24750 30960
rect 24980 31060 25040 31080
rect 24980 30900 24990 31060
rect 25030 30900 25040 31060
rect 23990 30880 24220 30900
rect 23990 30840 24150 30880
rect 24190 30840 24220 30880
rect 23990 30820 24220 30840
rect 24330 30880 24390 30900
rect 24330 30840 24340 30880
rect 24380 30840 24390 30880
rect 24330 30820 24390 30840
rect 24430 30880 24540 30900
rect 24430 30840 24490 30880
rect 24530 30840 24540 30880
rect 24430 30820 24540 30840
rect 24590 30880 24650 30900
rect 24590 30840 24600 30880
rect 24640 30840 24650 30880
rect 24590 30820 24650 30840
rect 24690 30880 24800 30900
rect 24690 30840 24740 30880
rect 24780 30840 24800 30880
rect 24690 30820 24800 30840
rect 24980 30840 25040 30900
rect 25090 31060 25150 31400
rect 25340 31320 25400 31550
rect 25340 31300 25480 31320
rect 25340 31260 25430 31300
rect 25470 31260 25480 31300
rect 25340 31240 25480 31260
rect 25090 30900 25100 31060
rect 25140 30900 25150 31060
rect 25090 30880 25150 30900
rect 25230 31060 25290 31080
rect 25230 30900 25240 31060
rect 25280 30900 25290 31060
rect 25230 30840 25290 30900
rect 25340 31060 25400 31240
rect 25340 30900 25350 31060
rect 25390 30900 25400 31060
rect 25340 30880 25400 30900
rect 23050 30390 23060 30550
rect 23100 30390 23110 30550
rect 23050 30370 23110 30390
rect 23160 30550 23220 30570
rect 23160 30390 23170 30550
rect 23210 30390 23220 30550
rect 23530 30550 23590 30570
rect 22690 30290 23120 30300
rect 22690 30250 22710 30290
rect 22750 30250 22890 30290
rect 22930 30250 23060 30290
rect 23100 30250 23120 30290
rect 22690 30240 23120 30250
rect 23160 30140 23220 30390
rect 23530 30390 23540 30550
rect 23580 30390 23590 30550
rect 23530 30140 23590 30390
rect 23640 30550 23700 30640
rect 23640 30390 23650 30550
rect 23690 30390 23700 30550
rect 23640 30370 23700 30390
rect 23990 30550 24050 30820
rect 24320 30760 24380 30780
rect 23990 30390 24000 30550
rect 24040 30390 24050 30550
rect 23990 30370 24050 30390
rect 24100 30550 24160 30570
rect 24100 30390 24110 30550
rect 24150 30390 24160 30550
rect 23630 30290 24060 30300
rect 23630 30250 23650 30290
rect 23690 30250 23830 30290
rect 23870 30250 24000 30290
rect 24040 30250 24060 30290
rect 23630 30240 24060 30250
rect 24100 30140 24160 30390
rect 24320 30400 24330 30760
rect 24370 30400 24380 30760
rect 24320 30140 24380 30400
rect 24430 30760 24490 30820
rect 24430 30400 24440 30760
rect 24480 30400 24490 30760
rect 24430 30380 24490 30400
rect 24580 30760 24640 30780
rect 24580 30400 24590 30760
rect 24630 30400 24640 30760
rect 24580 30140 24640 30400
rect 24690 30760 24750 30820
rect 24980 30800 25150 30840
rect 24690 30400 24700 30760
rect 24740 30400 24750 30760
rect 24950 30740 25050 30760
rect 24950 30680 24970 30740
rect 25030 30680 25050 30740
rect 24950 30660 25050 30680
rect 25090 30750 25150 30800
rect 25230 30790 25400 30840
rect 25090 30740 25300 30750
rect 25090 30700 25100 30740
rect 25140 30700 25240 30740
rect 25280 30700 25300 30740
rect 25090 30690 25300 30700
rect 24970 30590 25050 30600
rect 24970 30550 24990 30590
rect 25030 30550 25050 30590
rect 24970 30540 25050 30550
rect 24690 30380 24750 30400
rect 24980 30480 25040 30500
rect 24980 30320 24990 30480
rect 25030 30320 25040 30480
rect 24980 30140 25040 30320
rect 25090 30480 25150 30690
rect 25090 30320 25100 30480
rect 25140 30320 25150 30480
rect 25090 30300 25150 30320
rect 25340 30140 25400 30790
rect 11180 29910 11240 30120
rect 14830 30130 25680 30140
rect 14830 30060 14870 30130
rect 14930 30060 14970 30130
rect 15030 30060 15070 30130
rect 15130 30060 15170 30130
rect 15230 30060 15270 30130
rect 15330 30060 15370 30130
rect 15430 30060 15470 30130
rect 15530 30060 15570 30130
rect 15630 30060 15670 30130
rect 15730 30060 15780 30130
rect 15840 30060 15880 30130
rect 15940 30060 15990 30130
rect 16050 30060 16130 30130
rect 16190 30060 16270 30130
rect 16330 30060 16370 30130
rect 16430 30060 16470 30130
rect 16530 30060 16570 30130
rect 16630 30060 16670 30130
rect 16730 30060 16770 30130
rect 16830 30060 16870 30130
rect 16930 30060 16970 30130
rect 17030 30060 17070 30130
rect 17130 30060 17170 30130
rect 17230 30060 17270 30130
rect 17330 30060 17370 30130
rect 17430 30060 17470 30130
rect 17530 30060 17570 30130
rect 17630 30060 17670 30130
rect 17730 30060 17770 30130
rect 17830 30060 17870 30130
rect 17930 30060 17970 30130
rect 18030 30060 18070 30130
rect 18130 30060 18170 30130
rect 18230 30060 18270 30130
rect 18330 30060 18370 30130
rect 18430 30060 18470 30130
rect 18530 30060 18570 30130
rect 18630 30060 18670 30130
rect 18730 30060 18770 30130
rect 18830 30060 18870 30130
rect 18930 30060 18970 30130
rect 19030 30060 19070 30130
rect 19130 30060 19170 30130
rect 19230 30060 19270 30130
rect 19330 30060 19370 30130
rect 19430 30060 19470 30130
rect 19530 30060 19570 30130
rect 19630 30060 19670 30130
rect 19730 30060 19770 30130
rect 19830 30060 19870 30130
rect 19930 30060 19970 30130
rect 20030 30060 20070 30130
rect 20130 30060 20170 30130
rect 20230 30060 20270 30130
rect 20330 30060 20370 30130
rect 20430 30060 20470 30130
rect 20530 30060 20570 30130
rect 20630 30060 20670 30130
rect 20730 30060 20770 30130
rect 20830 30060 20870 30130
rect 20930 30060 20970 30130
rect 21030 30060 21070 30130
rect 21130 30060 21170 30130
rect 21230 30060 21270 30130
rect 21330 30060 21370 30130
rect 21430 30060 21470 30130
rect 21530 30060 21570 30130
rect 21630 30060 21670 30130
rect 21730 30060 21770 30130
rect 21830 30060 21870 30130
rect 21930 30060 21970 30130
rect 22030 30060 22070 30130
rect 22130 30060 22170 30130
rect 22230 30060 22270 30130
rect 22330 30060 22370 30130
rect 22430 30060 22470 30130
rect 22530 30060 22570 30130
rect 22630 30060 22670 30130
rect 22730 30060 22770 30130
rect 22830 30060 22870 30130
rect 22930 30060 22970 30130
rect 23030 30060 23070 30130
rect 23130 30060 23170 30130
rect 23230 30060 23270 30130
rect 23330 30060 23370 30130
rect 23430 30060 23470 30130
rect 23530 30060 23570 30130
rect 23630 30060 23670 30130
rect 23730 30060 23770 30130
rect 23830 30060 23870 30130
rect 23930 30060 23970 30130
rect 24030 30060 24070 30130
rect 24130 30060 24170 30130
rect 24230 30060 24270 30130
rect 24330 30060 24370 30130
rect 24430 30060 24470 30130
rect 24530 30060 24570 30130
rect 24630 30060 24670 30130
rect 24730 30060 24770 30130
rect 24830 30060 24870 30130
rect 24930 30060 24970 30130
rect 25030 30060 25070 30130
rect 25130 30060 25170 30130
rect 25230 30060 25270 30130
rect 25330 30060 25370 30130
rect 25430 30060 25470 30130
rect 25530 30060 25570 30130
rect 25630 30060 25680 30130
rect 14830 30050 25680 30060
rect 6400 29900 11240 29910
rect 6400 29840 6440 29900
rect 6500 29840 6540 29900
rect 6600 29840 6640 29900
rect 6700 29840 6740 29900
rect 6800 29840 6840 29900
rect 6900 29840 6940 29900
rect 7000 29840 7040 29900
rect 7100 29840 7140 29900
rect 7200 29840 7240 29900
rect 7300 29840 7340 29900
rect 7400 29840 7440 29900
rect 7500 29840 7540 29900
rect 7600 29840 7640 29900
rect 7700 29840 7740 29900
rect 7800 29840 7840 29900
rect 7900 29840 7940 29900
rect 8000 29840 8040 29900
rect 8100 29840 8140 29900
rect 8200 29840 8240 29900
rect 8300 29840 8340 29900
rect 8400 29840 8440 29900
rect 8500 29840 8540 29900
rect 8600 29840 8640 29900
rect 8700 29840 8740 29900
rect 8800 29840 8840 29900
rect 8900 29840 8940 29900
rect 9000 29840 9040 29900
rect 9100 29840 9140 29900
rect 9200 29840 9240 29900
rect 9300 29840 9340 29900
rect 9400 29840 9440 29900
rect 9500 29840 9540 29900
rect 9600 29840 9640 29900
rect 9700 29840 9740 29900
rect 9800 29840 9840 29900
rect 9900 29840 9940 29900
rect 10000 29840 10040 29900
rect 10100 29840 10140 29900
rect 10200 29840 10240 29900
rect 10300 29840 10340 29900
rect 10400 29840 10440 29900
rect 10500 29840 10540 29900
rect 10600 29840 10640 29900
rect 10700 29840 10740 29900
rect 10800 29840 10840 29900
rect 10900 29840 10940 29900
rect 11000 29840 11040 29900
rect 11100 29840 11140 29900
rect 11200 29840 11240 29900
rect 6400 29830 11240 29840
rect 6240 29510 6300 29530
rect 2170 29370 6310 29380
rect 2170 29310 2210 29370
rect 2270 29310 2310 29370
rect 2370 29310 2410 29370
rect 2470 29310 2510 29370
rect 2570 29310 2610 29370
rect 2670 29310 2710 29370
rect 2770 29310 2810 29370
rect 2870 29310 2910 29370
rect 2970 29310 3010 29370
rect 3070 29310 3110 29370
rect 3170 29310 3210 29370
rect 3270 29310 3310 29370
rect 3370 29310 3410 29370
rect 3470 29310 3510 29370
rect 3570 29310 3610 29370
rect 3670 29310 3710 29370
rect 3770 29310 3810 29370
rect 3870 29310 3910 29370
rect 3970 29310 4010 29370
rect 4070 29310 4110 29370
rect 4170 29310 4210 29370
rect 4270 29310 4310 29370
rect 4370 29310 4410 29370
rect 4470 29310 4510 29370
rect 4570 29310 4610 29370
rect 4670 29310 4710 29370
rect 4770 29310 4810 29370
rect 4870 29310 4910 29370
rect 4970 29310 5010 29370
rect 5070 29310 5110 29370
rect 5170 29310 5210 29370
rect 5270 29310 5310 29370
rect 5370 29310 5410 29370
rect 5470 29310 5510 29370
rect 5570 29310 5610 29370
rect 5670 29310 5710 29370
rect 5770 29310 5810 29370
rect 5870 29310 5910 29370
rect 5970 29310 6010 29370
rect 6070 29310 6110 29370
rect 6170 29310 6210 29370
rect 6270 29310 6310 29370
rect 2170 29300 6310 29310
rect 7320 26610 20640 26620
rect 7320 26570 7360 26610
rect 7400 26570 7440 26610
rect 7480 26570 7520 26610
rect 7560 26570 7600 26610
rect 7640 26570 7680 26610
rect 7720 26570 7760 26610
rect 7800 26570 7840 26610
rect 7880 26570 7920 26610
rect 7960 26570 8000 26610
rect 8040 26570 8080 26610
rect 8120 26570 8160 26610
rect 8200 26570 8240 26610
rect 8280 26570 8320 26610
rect 8360 26570 8400 26610
rect 8440 26570 8480 26610
rect 8520 26570 8560 26610
rect 8600 26570 8640 26610
rect 8680 26570 8720 26610
rect 8760 26570 8800 26610
rect 8840 26570 8880 26610
rect 8920 26570 8960 26610
rect 9000 26570 9040 26610
rect 9080 26570 9120 26610
rect 9160 26570 9200 26610
rect 9240 26570 9280 26610
rect 9320 26570 9360 26610
rect 9400 26570 9440 26610
rect 9480 26570 9520 26610
rect 9560 26570 9600 26610
rect 9640 26570 9680 26610
rect 9720 26570 9760 26610
rect 9800 26570 9840 26610
rect 9880 26570 9920 26610
rect 9960 26570 10000 26610
rect 10040 26570 10080 26610
rect 10120 26570 10160 26610
rect 10200 26570 10240 26610
rect 10280 26570 10320 26610
rect 10360 26570 10400 26610
rect 10440 26570 10480 26610
rect 10520 26570 10560 26610
rect 10600 26570 10640 26610
rect 10680 26570 10720 26610
rect 10760 26570 10800 26610
rect 10840 26570 10880 26610
rect 10920 26570 10960 26610
rect 11000 26570 11040 26610
rect 11080 26570 11120 26610
rect 11160 26570 11200 26610
rect 11240 26570 11280 26610
rect 11320 26570 11360 26610
rect 11400 26570 11440 26610
rect 11480 26570 11520 26610
rect 11560 26570 11600 26610
rect 11640 26570 11680 26610
rect 11720 26570 11760 26610
rect 11800 26570 11840 26610
rect 11880 26570 11920 26610
rect 11960 26570 12000 26610
rect 12040 26570 12080 26610
rect 12120 26570 12160 26610
rect 12200 26570 12240 26610
rect 12280 26570 12320 26610
rect 12360 26570 12400 26610
rect 12440 26570 12480 26610
rect 12520 26570 12560 26610
rect 12600 26570 12640 26610
rect 12680 26570 12720 26610
rect 12760 26570 12800 26610
rect 12840 26570 12880 26610
rect 12920 26570 12960 26610
rect 13000 26570 13040 26610
rect 13080 26570 13120 26610
rect 13160 26570 13200 26610
rect 13240 26570 13280 26610
rect 13320 26570 13360 26610
rect 13400 26570 13440 26610
rect 13480 26570 13520 26610
rect 13560 26570 13600 26610
rect 13640 26570 13680 26610
rect 13720 26570 13760 26610
rect 13800 26570 13840 26610
rect 13880 26570 13920 26610
rect 13960 26570 14000 26610
rect 14040 26570 14080 26610
rect 14120 26570 14160 26610
rect 14200 26570 14240 26610
rect 14280 26570 14320 26610
rect 14360 26570 14400 26610
rect 14440 26570 14480 26610
rect 14520 26570 14560 26610
rect 14600 26570 14640 26610
rect 14680 26570 14720 26610
rect 14760 26570 14800 26610
rect 14840 26570 14880 26610
rect 14920 26570 14960 26610
rect 15000 26570 15040 26610
rect 15080 26570 15120 26610
rect 15160 26570 15200 26610
rect 15240 26570 15280 26610
rect 15320 26570 15360 26610
rect 15400 26570 15440 26610
rect 15480 26570 15520 26610
rect 15560 26570 15600 26610
rect 15640 26570 15680 26610
rect 15720 26570 15760 26610
rect 15800 26570 15840 26610
rect 15880 26570 15920 26610
rect 15960 26570 16000 26610
rect 16040 26570 16080 26610
rect 16120 26570 16160 26610
rect 16200 26570 16240 26610
rect 16280 26570 16320 26610
rect 16360 26570 16400 26610
rect 16440 26570 16480 26610
rect 16520 26570 16560 26610
rect 16600 26570 16640 26610
rect 16680 26570 16720 26610
rect 16760 26570 16800 26610
rect 16840 26570 16880 26610
rect 16920 26570 16960 26610
rect 17000 26570 17040 26610
rect 17080 26570 17120 26610
rect 17160 26570 17200 26610
rect 17240 26570 17280 26610
rect 17320 26570 17360 26610
rect 17400 26570 17440 26610
rect 17480 26570 17520 26610
rect 17560 26570 17600 26610
rect 17640 26570 17680 26610
rect 17720 26570 17760 26610
rect 17800 26570 17840 26610
rect 17880 26570 17920 26610
rect 17960 26570 18000 26610
rect 18040 26570 18080 26610
rect 18120 26570 18160 26610
rect 18200 26570 18240 26610
rect 18280 26570 18320 26610
rect 18360 26570 18400 26610
rect 18440 26570 18480 26610
rect 18520 26570 18560 26610
rect 18600 26570 18640 26610
rect 18680 26570 18720 26610
rect 18760 26570 18800 26610
rect 18840 26570 18880 26610
rect 18920 26570 18960 26610
rect 19000 26570 19040 26610
rect 19080 26570 19120 26610
rect 19160 26570 19200 26610
rect 19240 26570 19280 26610
rect 19320 26570 19360 26610
rect 19400 26570 19440 26610
rect 19480 26570 19520 26610
rect 19560 26570 19600 26610
rect 19640 26570 19680 26610
rect 19720 26570 19760 26610
rect 19800 26570 19840 26610
rect 19880 26570 19920 26610
rect 19960 26570 20000 26610
rect 20040 26570 20080 26610
rect 20120 26570 20160 26610
rect 20200 26570 20240 26610
rect 20280 26570 20320 26610
rect 20360 26570 20400 26610
rect 20440 26570 20480 26610
rect 20520 26570 20560 26610
rect 20600 26570 20640 26610
rect 7320 26560 20640 26570
rect 7320 26470 7380 26560
rect 7320 26010 7330 26470
rect 7370 26010 7380 26470
rect 7320 25990 7380 26010
rect 7430 26470 7490 26490
rect 7430 26010 7440 26470
rect 7480 26010 7490 26470
rect 6280 25560 7160 25580
rect 6280 25500 6300 25560
rect 6360 25500 7080 25560
rect 7140 25500 7160 25560
rect 6280 25480 7160 25500
rect 7270 25190 7390 25210
rect 7270 25130 7290 25190
rect 7350 25130 7390 25190
rect 7270 25110 7390 25130
rect 7430 24790 7490 26010
rect 7540 26470 7600 26560
rect 7540 26010 7550 26470
rect 7590 26010 7600 26470
rect 7540 25990 7600 26010
rect 7850 26470 7910 26560
rect 7850 26010 7860 26470
rect 7900 26010 7910 26470
rect 7850 25990 7910 26010
rect 7960 26470 8020 26490
rect 7960 26010 7970 26470
rect 8010 26010 8020 26470
rect 7800 25560 7920 25580
rect 7800 25500 7820 25560
rect 7880 25500 7920 25560
rect 7800 25480 7920 25500
rect 7960 24860 8020 26010
rect 8070 26470 8130 26560
rect 8070 26010 8080 26470
rect 8120 26010 8130 26470
rect 8070 25990 8130 26010
rect 8480 26480 8540 26560
rect 8480 26020 8490 26480
rect 8530 26020 8540 26480
rect 8480 26000 8540 26020
rect 8610 26480 8670 26500
rect 8610 26020 8620 26480
rect 8660 26020 8670 26480
rect 8610 24960 8670 26020
rect 8740 26480 8800 26560
rect 8740 26020 8750 26480
rect 8790 26020 8800 26480
rect 8740 26000 8800 26020
rect 8860 26480 8920 26560
rect 8860 26020 8870 26480
rect 8910 26020 8920 26480
rect 8860 26000 8920 26020
rect 8970 26480 9030 26500
rect 8970 26020 8980 26480
rect 9020 26020 9030 26480
rect 8970 24960 9030 26020
rect 9220 26480 9280 26560
rect 9220 26020 9230 26480
rect 9270 26020 9280 26480
rect 9220 26000 9280 26020
rect 9330 26480 9390 26500
rect 9330 26020 9340 26480
rect 9380 26020 9390 26480
rect 8480 24940 8550 24960
rect 8480 24900 8500 24940
rect 8540 24900 8550 24940
rect 8610 24940 8930 24960
rect 8610 24920 8800 24940
rect 8480 24880 8550 24900
rect 8740 24900 8800 24920
rect 8840 24900 8880 24940
rect 8920 24900 8930 24940
rect 8740 24880 8930 24900
rect 8970 24950 9160 24960
rect 8970 24890 8990 24950
rect 9050 24890 9160 24950
rect 9200 24950 9290 24960
rect 9200 24910 9220 24950
rect 9260 24910 9290 24950
rect 9200 24900 9290 24910
rect 8970 24880 9160 24890
rect 8060 24870 8160 24880
rect 8060 24860 8080 24870
rect 7960 24800 8080 24860
rect 8140 24800 8160 24870
rect 8630 24860 8700 24880
rect 8630 24820 8650 24860
rect 8690 24820 8700 24860
rect 8630 24800 8700 24820
rect 7430 24770 7650 24790
rect 7430 24710 7570 24770
rect 7630 24710 7650 24770
rect 7430 24690 7650 24710
rect 7320 24550 7380 24570
rect 7320 24390 7330 24550
rect 7370 24390 7380 24550
rect 7320 24300 7380 24390
rect 7430 24550 7490 24690
rect 7430 24390 7440 24550
rect 7480 24390 7490 24550
rect 7430 24370 7490 24390
rect 7540 24550 7600 24570
rect 7540 24390 7550 24550
rect 7590 24390 7600 24550
rect 7540 24300 7600 24390
rect 7850 24550 7910 24570
rect 7850 24390 7860 24550
rect 7900 24390 7910 24550
rect 7850 24300 7910 24390
rect 7960 24550 8020 24800
rect 8060 24790 8160 24800
rect 8180 24730 8280 24750
rect 8180 24670 8200 24730
rect 8260 24670 8280 24730
rect 8180 24650 8280 24670
rect 8480 24740 8540 24760
rect 7960 24390 7970 24550
rect 8010 24390 8020 24550
rect 7960 24370 8020 24390
rect 8070 24550 8130 24570
rect 8070 24390 8080 24550
rect 8120 24390 8130 24550
rect 8070 24300 8130 24390
rect 8480 24380 8490 24740
rect 8530 24380 8540 24740
rect 8480 24300 8540 24380
rect 8610 24740 8670 24760
rect 8610 24380 8620 24740
rect 8660 24380 8670 24740
rect 8610 24360 8670 24380
rect 8740 24740 8800 24880
rect 8740 24380 8750 24740
rect 8790 24380 8800 24740
rect 8740 24360 8800 24380
rect 8860 24810 8920 24830
rect 8860 24650 8870 24810
rect 8910 24650 8920 24810
rect 8860 24300 8920 24650
rect 8970 24810 9030 24880
rect 8970 24650 8980 24810
rect 9020 24650 9030 24810
rect 8970 24630 9030 24650
rect 9090 24630 9160 24880
rect 9330 24840 9390 26020
rect 9440 26480 9500 26560
rect 9440 26020 9450 26480
rect 9490 26020 9500 26480
rect 9440 26000 9500 26020
rect 9670 26480 9730 26560
rect 9670 26020 9680 26480
rect 9720 26020 9730 26480
rect 9670 26000 9730 26020
rect 9800 26480 9860 26500
rect 9800 26020 9810 26480
rect 9850 26020 9860 26480
rect 9660 25950 9740 25960
rect 9660 25910 9680 25950
rect 9720 25910 9740 25950
rect 9660 25900 9740 25910
rect 9660 25060 9740 25070
rect 9660 25020 9680 25060
rect 9720 25020 9740 25060
rect 9660 25010 9740 25020
rect 9800 24960 9860 26020
rect 9930 26480 9990 26560
rect 9930 26020 9940 26480
rect 9980 26020 9990 26480
rect 9930 26000 9990 26020
rect 10160 26480 10220 26560
rect 10160 26020 10170 26480
rect 10210 26020 10220 26480
rect 10160 26000 10220 26020
rect 10270 26480 10330 26500
rect 10270 26020 10280 26480
rect 10320 26020 10330 26480
rect 9920 25950 10000 25960
rect 9920 25910 9940 25950
rect 9980 25910 10000 25950
rect 9920 25900 10000 25910
rect 9920 25060 10000 25070
rect 9920 25020 9940 25060
rect 9980 25020 10000 25060
rect 9920 25010 10000 25020
rect 10270 24960 10330 26020
rect 10380 26480 10440 26560
rect 10380 26020 10390 26480
rect 10430 26020 10440 26480
rect 10380 26000 10440 26020
rect 10660 26480 10720 26560
rect 10660 26020 10670 26480
rect 10710 26020 10720 26480
rect 10660 26000 10720 26020
rect 10790 26480 10850 26500
rect 10790 26020 10800 26480
rect 10840 26020 10850 26480
rect 10650 25950 10730 25960
rect 10650 25910 10670 25950
rect 10710 25910 10730 25950
rect 10650 25900 10730 25910
rect 10650 25060 10730 25070
rect 10650 25020 10670 25060
rect 10710 25020 10730 25060
rect 10650 25010 10730 25020
rect 10790 24960 10850 26020
rect 10920 26480 10980 26560
rect 10920 26020 10930 26480
rect 10970 26020 10980 26480
rect 10920 26000 10980 26020
rect 11150 26480 11210 26560
rect 11150 26020 11160 26480
rect 11200 26020 11210 26480
rect 11150 26000 11210 26020
rect 11260 26480 11320 26500
rect 11260 26020 11270 26480
rect 11310 26020 11320 26480
rect 10910 25950 10990 25960
rect 10910 25910 10930 25950
rect 10970 25910 10990 25950
rect 10910 25900 10990 25910
rect 10910 25060 10990 25070
rect 10910 25020 10930 25060
rect 10970 25020 10990 25060
rect 10910 25010 10990 25020
rect 11260 24960 11320 26020
rect 11370 26480 11430 26560
rect 11370 26020 11380 26480
rect 11420 26020 11430 26480
rect 11370 26000 11430 26020
rect 11660 26480 11720 26560
rect 11660 26020 11670 26480
rect 11710 26020 11720 26480
rect 11660 26000 11720 26020
rect 11790 26480 11850 26500
rect 11790 26020 11800 26480
rect 11840 26020 11850 26480
rect 11650 25950 11730 25960
rect 11650 25910 11670 25950
rect 11710 25910 11730 25950
rect 11650 25900 11730 25910
rect 11650 25060 11730 25070
rect 11650 25020 11670 25060
rect 11710 25020 11730 25060
rect 11650 25010 11730 25020
rect 11790 24960 11850 26020
rect 11920 26480 11980 26560
rect 11920 26020 11930 26480
rect 11970 26020 11980 26480
rect 11920 26000 11980 26020
rect 12150 26480 12210 26560
rect 12150 26020 12160 26480
rect 12200 26020 12210 26480
rect 12150 26000 12210 26020
rect 12260 26480 12320 26500
rect 12260 26020 12270 26480
rect 12310 26020 12320 26480
rect 11910 25950 11990 25960
rect 11910 25910 11930 25950
rect 11970 25910 11990 25950
rect 11910 25900 11990 25910
rect 11910 25060 11990 25070
rect 11910 25020 11930 25060
rect 11970 25020 11990 25060
rect 11910 25010 11990 25020
rect 12260 24960 12320 26020
rect 12370 26480 12430 26560
rect 12370 26020 12380 26480
rect 12420 26020 12430 26480
rect 12370 26000 12430 26020
rect 12530 26480 12590 26560
rect 12530 26020 12540 26480
rect 12580 26020 12590 26480
rect 12530 26000 12590 26020
rect 12640 26480 12700 26500
rect 12640 26020 12650 26480
rect 12690 26020 12700 26480
rect 12640 24960 12700 26020
rect 12750 26480 12810 26560
rect 12750 26020 12760 26480
rect 12800 26020 12810 26480
rect 12750 26000 12810 26020
rect 12880 26480 12940 26560
rect 12880 26020 12890 26480
rect 12930 26020 12940 26480
rect 12880 26000 12940 26020
rect 12990 26480 13050 26500
rect 12990 26020 13000 26480
rect 13040 26020 13050 26480
rect 9570 24940 9630 24960
rect 9570 24900 9580 24940
rect 9620 24900 9630 24940
rect 9800 24950 10230 24960
rect 9800 24910 10080 24950
rect 10120 24910 10160 24950
rect 10200 24910 10230 24950
rect 9800 24900 10230 24910
rect 10270 24950 10510 24960
rect 10270 24910 10460 24950
rect 10500 24910 10510 24950
rect 10270 24900 10510 24910
rect 10560 24940 10620 24960
rect 10560 24900 10570 24940
rect 10610 24900 10620 24940
rect 10790 24950 11220 24960
rect 10790 24910 11070 24950
rect 11110 24910 11150 24950
rect 11190 24910 11220 24950
rect 10790 24900 11220 24910
rect 11260 24950 11500 24960
rect 11260 24910 11450 24950
rect 11490 24910 11500 24950
rect 11260 24900 11500 24910
rect 11560 24940 11620 24960
rect 11560 24900 11570 24940
rect 11610 24900 11620 24940
rect 11790 24950 12220 24960
rect 11790 24910 12070 24950
rect 12110 24910 12150 24950
rect 12190 24910 12220 24950
rect 11790 24900 12220 24910
rect 12260 24950 12600 24960
rect 12260 24910 12450 24950
rect 12490 24910 12530 24950
rect 12570 24910 12600 24950
rect 12260 24900 12600 24910
rect 12640 24940 12950 24960
rect 12640 24900 12820 24940
rect 12860 24900 12900 24940
rect 12940 24900 12950 24940
rect 9570 24880 9630 24900
rect 9830 24840 9890 24860
rect 9330 24800 9840 24840
rect 9880 24800 9890 24840
rect 9080 24610 9170 24630
rect 9080 24560 9100 24610
rect 9150 24560 9170 24610
rect 9080 24540 9170 24560
rect 9220 24540 9280 24560
rect 9220 24380 9230 24540
rect 9270 24380 9280 24540
rect 9220 24300 9280 24380
rect 9330 24540 9390 24800
rect 9830 24780 9890 24800
rect 9670 24740 9730 24760
rect 9330 24380 9340 24540
rect 9380 24380 9390 24540
rect 9330 24360 9390 24380
rect 9440 24540 9500 24560
rect 9440 24380 9450 24540
rect 9490 24380 9500 24540
rect 9440 24300 9500 24380
rect 9670 24380 9680 24740
rect 9720 24380 9730 24740
rect 9670 24300 9730 24380
rect 9930 24740 9990 24900
rect 9930 24380 9940 24740
rect 9980 24380 9990 24740
rect 9930 24360 9990 24380
rect 10160 24540 10220 24560
rect 10160 24380 10170 24540
rect 10210 24380 10220 24540
rect 10160 24300 10220 24380
rect 10270 24540 10330 24900
rect 10560 24880 10620 24900
rect 10820 24840 10880 24860
rect 10820 24800 10830 24840
rect 10870 24800 10880 24840
rect 10820 24780 10880 24800
rect 10660 24740 10720 24760
rect 10270 24380 10280 24540
rect 10320 24380 10330 24540
rect 10270 24360 10330 24380
rect 10380 24540 10440 24560
rect 10380 24380 10390 24540
rect 10430 24380 10440 24540
rect 10380 24300 10440 24380
rect 10660 24380 10670 24740
rect 10710 24380 10720 24740
rect 10660 24300 10720 24380
rect 10920 24740 10980 24900
rect 10920 24380 10930 24740
rect 10970 24380 10980 24740
rect 10920 24360 10980 24380
rect 11150 24540 11210 24560
rect 11150 24380 11160 24540
rect 11200 24380 11210 24540
rect 11150 24300 11210 24380
rect 11260 24540 11320 24900
rect 11560 24880 11620 24900
rect 11820 24840 11880 24860
rect 11820 24800 11830 24840
rect 11870 24800 11880 24840
rect 11820 24780 11880 24800
rect 11660 24740 11720 24760
rect 11260 24380 11270 24540
rect 11310 24380 11320 24540
rect 11260 24360 11320 24380
rect 11370 24540 11430 24560
rect 11370 24380 11380 24540
rect 11420 24380 11430 24540
rect 11370 24300 11430 24380
rect 11660 24380 11670 24740
rect 11710 24380 11720 24740
rect 11660 24300 11720 24380
rect 11920 24740 11980 24900
rect 11920 24380 11930 24740
rect 11970 24380 11980 24740
rect 11920 24360 11980 24380
rect 12150 24540 12210 24560
rect 12150 24380 12160 24540
rect 12200 24380 12210 24540
rect 12150 24300 12210 24380
rect 12260 24540 12320 24900
rect 12640 24880 12950 24900
rect 12990 24940 13050 26020
rect 13110 26480 13170 26500
rect 13110 26020 13120 26480
rect 13160 26020 13170 26480
rect 13110 26000 13170 26020
rect 13220 26480 13280 26560
rect 13220 26020 13230 26480
rect 13270 26020 13280 26480
rect 13220 26000 13280 26020
rect 13330 26480 13390 26500
rect 13330 26020 13340 26480
rect 13380 26020 13390 26480
rect 13210 25930 13290 25940
rect 13210 25890 13230 25930
rect 13270 25890 13290 25930
rect 13210 25880 13290 25890
rect 13210 25040 13290 25050
rect 13210 25000 13230 25040
rect 13270 25000 13290 25040
rect 13210 24990 13290 25000
rect 12990 24900 13000 24940
rect 13040 24900 13050 24940
rect 12260 24380 12270 24540
rect 12310 24380 12320 24540
rect 12260 24360 12320 24380
rect 12370 24540 12430 24560
rect 12370 24380 12380 24540
rect 12420 24380 12430 24540
rect 12370 24300 12430 24380
rect 12530 24540 12590 24560
rect 12530 24380 12540 24540
rect 12580 24380 12590 24540
rect 12530 24300 12590 24380
rect 12640 24540 12700 24880
rect 12880 24820 12940 24840
rect 12880 24660 12890 24820
rect 12930 24660 12940 24820
rect 12640 24380 12650 24540
rect 12690 24380 12700 24540
rect 12640 24360 12700 24380
rect 12750 24540 12810 24560
rect 12750 24380 12760 24540
rect 12800 24380 12810 24540
rect 12750 24300 12810 24380
rect 12880 24300 12940 24660
rect 12990 24820 13050 24900
rect 13120 24940 13180 24960
rect 13120 24900 13130 24940
rect 13170 24900 13180 24940
rect 13120 24880 13180 24900
rect 13330 24940 13390 26020
rect 13450 26480 13510 26500
rect 13450 26020 13460 26480
rect 13500 26020 13510 26480
rect 13450 26000 13510 26020
rect 13560 26480 13620 26560
rect 13560 26020 13570 26480
rect 13610 26020 13620 26480
rect 13560 26000 13620 26020
rect 13670 26480 13730 26500
rect 13670 26020 13680 26480
rect 13720 26020 13730 26480
rect 13670 26000 13730 26020
rect 13780 26480 13840 26560
rect 13780 26020 13790 26480
rect 13830 26020 13840 26480
rect 13780 26000 13840 26020
rect 13890 26480 13950 26500
rect 13890 26020 13900 26480
rect 13940 26020 13950 26480
rect 13550 25930 13630 25940
rect 13550 25890 13570 25930
rect 13610 25890 13630 25930
rect 13550 25880 13630 25890
rect 13770 25930 13850 25940
rect 13770 25890 13790 25930
rect 13830 25890 13850 25930
rect 13770 25880 13850 25890
rect 13550 25040 13630 25050
rect 13550 25000 13570 25040
rect 13610 25000 13630 25040
rect 13550 24990 13630 25000
rect 13770 25040 13850 25050
rect 13770 25000 13790 25040
rect 13830 25000 13850 25040
rect 13770 24990 13850 25000
rect 13330 24900 13340 24940
rect 13380 24900 13390 24940
rect 12990 24660 13000 24820
rect 13040 24660 13050 24820
rect 12990 24640 13050 24660
rect 13110 24820 13170 24840
rect 13110 24660 13120 24820
rect 13160 24660 13170 24820
rect 13110 24640 13170 24660
rect 13220 24820 13280 24840
rect 13220 24660 13230 24820
rect 13270 24660 13280 24820
rect 13220 24300 13280 24660
rect 13330 24820 13390 24900
rect 13460 24940 13520 24960
rect 13460 24900 13470 24940
rect 13510 24900 13520 24940
rect 13460 24880 13520 24900
rect 13890 24940 13950 26020
rect 14010 26480 14070 26500
rect 14010 26020 14020 26480
rect 14060 26020 14070 26480
rect 14010 26000 14070 26020
rect 14120 26480 14180 26560
rect 14120 26020 14130 26480
rect 14170 26020 14180 26480
rect 14120 26000 14180 26020
rect 14230 26480 14290 26500
rect 14230 26020 14240 26480
rect 14280 26020 14290 26480
rect 14230 26000 14290 26020
rect 14340 26480 14400 26560
rect 14340 26020 14350 26480
rect 14390 26020 14400 26480
rect 14340 26000 14400 26020
rect 14450 26480 14510 26500
rect 14450 26020 14460 26480
rect 14500 26020 14510 26480
rect 14450 26000 14510 26020
rect 14560 26480 14620 26560
rect 14560 26020 14570 26480
rect 14610 26020 14620 26480
rect 14560 26000 14620 26020
rect 14670 26480 14730 26500
rect 14670 26020 14680 26480
rect 14720 26020 14730 26480
rect 14670 26000 14730 26020
rect 14780 26480 14840 26560
rect 14780 26020 14790 26480
rect 14830 26020 14840 26480
rect 14780 26000 14840 26020
rect 14890 26480 14950 26500
rect 14890 26020 14900 26480
rect 14940 26020 14950 26480
rect 14110 25950 14190 25960
rect 14110 25910 14130 25950
rect 14170 25910 14190 25950
rect 14110 25900 14190 25910
rect 14330 25950 14410 25960
rect 14330 25910 14350 25950
rect 14390 25910 14410 25950
rect 14330 25900 14410 25910
rect 14550 25950 14630 25960
rect 14550 25910 14570 25950
rect 14610 25910 14630 25950
rect 14550 25900 14630 25910
rect 14770 25950 14850 25960
rect 14770 25910 14790 25950
rect 14830 25910 14850 25950
rect 14770 25900 14850 25910
rect 14110 25060 14190 25070
rect 14110 25020 14130 25060
rect 14170 25020 14190 25060
rect 14110 25010 14190 25020
rect 14330 25060 14410 25070
rect 14330 25020 14350 25060
rect 14390 25020 14410 25060
rect 14330 25010 14410 25020
rect 14550 25060 14630 25070
rect 14550 25020 14570 25060
rect 14610 25020 14630 25060
rect 14550 25010 14630 25020
rect 14770 25060 14850 25070
rect 14770 25020 14790 25060
rect 14830 25020 14850 25060
rect 14770 25010 14850 25020
rect 13890 24900 13900 24940
rect 13940 24900 13950 24940
rect 13330 24660 13340 24820
rect 13380 24660 13390 24820
rect 13330 24640 13390 24660
rect 13450 24820 13510 24840
rect 13450 24660 13460 24820
rect 13500 24660 13510 24820
rect 13450 24640 13510 24660
rect 13560 24820 13620 24840
rect 13560 24660 13570 24820
rect 13610 24660 13620 24820
rect 13560 24300 13620 24660
rect 13670 24820 13730 24840
rect 13670 24660 13680 24820
rect 13720 24660 13730 24820
rect 13670 24640 13730 24660
rect 13780 24820 13840 24840
rect 13780 24660 13790 24820
rect 13830 24660 13840 24820
rect 13780 24300 13840 24660
rect 13890 24820 13950 24900
rect 14020 24940 14080 24960
rect 14020 24900 14030 24940
rect 14070 24900 14080 24940
rect 14020 24880 14080 24900
rect 14890 24940 14950 26020
rect 15070 26480 15130 26500
rect 15070 26020 15080 26480
rect 15120 26020 15130 26480
rect 15070 26000 15130 26020
rect 15180 26480 15240 26560
rect 15180 26020 15190 26480
rect 15230 26020 15240 26480
rect 15180 26000 15240 26020
rect 15290 26480 15350 26500
rect 15290 26020 15300 26480
rect 15340 26020 15350 26480
rect 15290 26000 15350 26020
rect 15400 26480 15460 26560
rect 15400 26020 15410 26480
rect 15450 26020 15460 26480
rect 15400 26000 15460 26020
rect 15510 26480 15570 26500
rect 15510 26020 15520 26480
rect 15560 26020 15570 26480
rect 15510 26000 15570 26020
rect 15620 26480 15680 26560
rect 15620 26020 15630 26480
rect 15670 26020 15680 26480
rect 15620 26000 15680 26020
rect 15730 26480 15790 26500
rect 15730 26020 15740 26480
rect 15780 26020 15790 26480
rect 15730 26000 15790 26020
rect 15840 26480 15900 26560
rect 15840 26020 15850 26480
rect 15890 26020 15900 26480
rect 15840 26000 15900 26020
rect 15950 26480 16010 26500
rect 15950 26020 15960 26480
rect 16000 26020 16010 26480
rect 15950 26000 16010 26020
rect 16060 26480 16120 26560
rect 16060 26020 16070 26480
rect 16110 26020 16120 26480
rect 16060 26000 16120 26020
rect 16170 26480 16230 26500
rect 16170 26020 16180 26480
rect 16220 26020 16230 26480
rect 16170 26000 16230 26020
rect 16280 26480 16340 26560
rect 16280 26020 16290 26480
rect 16330 26020 16340 26480
rect 16280 26000 16340 26020
rect 16390 26480 16450 26500
rect 16390 26020 16400 26480
rect 16440 26020 16450 26480
rect 16390 26000 16450 26020
rect 16500 26480 16560 26560
rect 16500 26020 16510 26480
rect 16550 26020 16560 26480
rect 16500 26000 16560 26020
rect 16610 26480 16670 26500
rect 16610 26020 16620 26480
rect 16660 26020 16670 26480
rect 16610 26000 16670 26020
rect 16720 26480 16780 26560
rect 16720 26020 16730 26480
rect 16770 26020 16780 26480
rect 16720 26000 16780 26020
rect 16830 26480 16890 26500
rect 16830 26020 16840 26480
rect 16880 26020 16890 26480
rect 15170 25950 15250 25960
rect 15170 25910 15190 25950
rect 15230 25910 15250 25950
rect 15170 25900 15250 25910
rect 15390 25950 15470 25960
rect 15390 25910 15410 25950
rect 15450 25910 15470 25950
rect 15390 25900 15470 25910
rect 15610 25950 15690 25960
rect 15610 25910 15630 25950
rect 15670 25910 15690 25950
rect 15610 25900 15690 25910
rect 15830 25950 15910 25960
rect 15830 25910 15850 25950
rect 15890 25910 15910 25950
rect 15830 25900 15910 25910
rect 16050 25950 16130 25960
rect 16050 25910 16070 25950
rect 16110 25910 16130 25950
rect 16050 25900 16130 25910
rect 16270 25950 16350 25960
rect 16270 25910 16290 25950
rect 16330 25910 16350 25950
rect 16270 25900 16350 25910
rect 16490 25950 16570 25960
rect 16490 25910 16510 25950
rect 16550 25910 16570 25950
rect 16490 25900 16570 25910
rect 16710 25950 16790 25960
rect 16710 25910 16730 25950
rect 16770 25910 16790 25950
rect 16710 25900 16790 25910
rect 15170 25060 15250 25070
rect 15170 25020 15190 25060
rect 15230 25020 15250 25060
rect 15170 25010 15250 25020
rect 15390 25060 15470 25070
rect 15390 25020 15410 25060
rect 15450 25020 15470 25060
rect 15390 25010 15470 25020
rect 15610 25060 15690 25070
rect 15610 25020 15630 25060
rect 15670 25020 15690 25060
rect 15610 25010 15690 25020
rect 15830 25060 15910 25070
rect 15830 25020 15850 25060
rect 15890 25020 15910 25060
rect 15830 25010 15910 25020
rect 16050 25060 16130 25070
rect 16050 25020 16070 25060
rect 16110 25020 16130 25060
rect 16050 25010 16130 25020
rect 16270 25060 16350 25070
rect 16270 25020 16290 25060
rect 16330 25020 16350 25060
rect 16270 25010 16350 25020
rect 16490 25060 16570 25070
rect 16490 25020 16510 25060
rect 16550 25020 16570 25060
rect 16490 25010 16570 25020
rect 16710 25060 16790 25070
rect 16710 25020 16730 25060
rect 16770 25020 16790 25060
rect 16710 25010 16790 25020
rect 14890 24900 14900 24940
rect 14940 24900 14950 24940
rect 13890 24660 13900 24820
rect 13940 24660 13950 24820
rect 13890 24640 13950 24660
rect 14010 24820 14070 24840
rect 14010 24660 14020 24820
rect 14060 24660 14070 24820
rect 14010 24640 14070 24660
rect 14120 24820 14180 24840
rect 14120 24660 14130 24820
rect 14170 24660 14180 24820
rect 14120 24300 14180 24660
rect 14230 24820 14290 24840
rect 14230 24660 14240 24820
rect 14280 24660 14290 24820
rect 14230 24640 14290 24660
rect 14340 24820 14400 24840
rect 14340 24660 14350 24820
rect 14390 24660 14400 24820
rect 14340 24300 14400 24660
rect 14450 24820 14510 24840
rect 14450 24660 14460 24820
rect 14500 24660 14510 24820
rect 14450 24640 14510 24660
rect 14560 24820 14620 24840
rect 14560 24660 14570 24820
rect 14610 24660 14620 24820
rect 14560 24300 14620 24660
rect 14670 24820 14730 24840
rect 14670 24660 14680 24820
rect 14720 24660 14730 24820
rect 14670 24640 14730 24660
rect 14780 24820 14840 24840
rect 14780 24660 14790 24820
rect 14830 24660 14840 24820
rect 14780 24300 14840 24660
rect 14890 24820 14950 24900
rect 15080 24940 15140 24960
rect 15080 24900 15090 24940
rect 15130 24900 15140 24940
rect 15080 24880 15140 24900
rect 16830 24950 16890 26020
rect 17020 26480 17080 26500
rect 17020 26020 17030 26480
rect 17070 26020 17080 26480
rect 17020 26000 17080 26020
rect 17130 26480 17190 26560
rect 17130 26020 17140 26480
rect 17180 26020 17190 26480
rect 17130 26000 17190 26020
rect 17240 26480 17300 26500
rect 17240 26020 17250 26480
rect 17290 26020 17300 26480
rect 17240 26000 17300 26020
rect 17350 26480 17410 26560
rect 17350 26020 17360 26480
rect 17400 26020 17410 26480
rect 17350 26000 17410 26020
rect 17460 26480 17520 26500
rect 17460 26020 17470 26480
rect 17510 26020 17520 26480
rect 17460 26000 17520 26020
rect 17570 26480 17630 26560
rect 17570 26020 17580 26480
rect 17620 26020 17630 26480
rect 17570 26000 17630 26020
rect 17680 26480 17740 26500
rect 17680 26020 17690 26480
rect 17730 26020 17740 26480
rect 17680 26000 17740 26020
rect 17790 26480 17850 26560
rect 17790 26020 17800 26480
rect 17840 26020 17850 26480
rect 17790 26000 17850 26020
rect 17900 26480 17960 26500
rect 17900 26020 17910 26480
rect 17950 26020 17960 26480
rect 17900 26000 17960 26020
rect 18010 26480 18070 26560
rect 18010 26020 18020 26480
rect 18060 26020 18070 26480
rect 18010 26000 18070 26020
rect 18120 26480 18180 26500
rect 18120 26020 18130 26480
rect 18170 26020 18180 26480
rect 18120 26000 18180 26020
rect 18230 26480 18290 26560
rect 18230 26020 18240 26480
rect 18280 26020 18290 26480
rect 18230 26000 18290 26020
rect 18340 26480 18400 26500
rect 18340 26020 18350 26480
rect 18390 26020 18400 26480
rect 18340 26000 18400 26020
rect 18450 26480 18510 26560
rect 18450 26020 18460 26480
rect 18500 26020 18510 26480
rect 18450 26000 18510 26020
rect 18560 26480 18620 26500
rect 18560 26020 18570 26480
rect 18610 26020 18620 26480
rect 18560 26000 18620 26020
rect 18670 26480 18730 26560
rect 18670 26020 18680 26480
rect 18720 26020 18730 26480
rect 18670 26000 18730 26020
rect 18780 26480 18840 26500
rect 18780 26020 18790 26480
rect 18830 26020 18840 26480
rect 18780 26000 18840 26020
rect 18890 26480 18950 26560
rect 18890 26020 18900 26480
rect 18940 26020 18950 26480
rect 18890 26000 18950 26020
rect 19000 26480 19060 26500
rect 19000 26020 19010 26480
rect 19050 26020 19060 26480
rect 19000 26000 19060 26020
rect 19110 26480 19170 26560
rect 19110 26020 19120 26480
rect 19160 26020 19170 26480
rect 19110 26000 19170 26020
rect 19220 26480 19280 26500
rect 19220 26020 19230 26480
rect 19270 26020 19280 26480
rect 19220 26000 19280 26020
rect 19330 26480 19390 26560
rect 19330 26020 19340 26480
rect 19380 26020 19390 26480
rect 19330 26000 19390 26020
rect 19440 26480 19500 26500
rect 19440 26020 19450 26480
rect 19490 26020 19500 26480
rect 19440 26000 19500 26020
rect 19550 26480 19610 26560
rect 19550 26020 19560 26480
rect 19600 26020 19610 26480
rect 19550 26000 19610 26020
rect 19660 26480 19720 26500
rect 19660 26020 19670 26480
rect 19710 26020 19720 26480
rect 19660 26000 19720 26020
rect 19770 26480 19830 26560
rect 19770 26020 19780 26480
rect 19820 26020 19830 26480
rect 19770 26000 19830 26020
rect 19880 26480 19940 26500
rect 19880 26020 19890 26480
rect 19930 26020 19940 26480
rect 19880 26000 19940 26020
rect 19990 26480 20050 26560
rect 19990 26020 20000 26480
rect 20040 26020 20050 26480
rect 19990 26000 20050 26020
rect 20100 26480 20160 26500
rect 20100 26020 20110 26480
rect 20150 26020 20160 26480
rect 20100 26000 20160 26020
rect 20210 26480 20270 26560
rect 20210 26020 20220 26480
rect 20260 26020 20270 26480
rect 20210 26000 20270 26020
rect 20320 26480 20380 26500
rect 20320 26020 20330 26480
rect 20370 26020 20380 26480
rect 20320 26000 20380 26020
rect 20430 26480 20490 26560
rect 20430 26020 20440 26480
rect 20480 26020 20490 26480
rect 20430 26000 20490 26020
rect 20540 26480 20600 26500
rect 20540 26020 20550 26480
rect 20590 26020 20600 26480
rect 17120 25950 17200 25960
rect 17120 25910 17140 25950
rect 17180 25910 17200 25950
rect 17120 25900 17200 25910
rect 17340 25950 17420 25960
rect 17340 25910 17360 25950
rect 17400 25910 17420 25950
rect 17340 25900 17420 25910
rect 17560 25950 17640 25960
rect 17560 25910 17580 25950
rect 17620 25910 17640 25950
rect 17560 25900 17640 25910
rect 17780 25950 17860 25960
rect 17780 25910 17800 25950
rect 17840 25910 17860 25950
rect 17780 25900 17860 25910
rect 18000 25950 18080 25960
rect 18000 25910 18020 25950
rect 18060 25910 18080 25950
rect 18000 25900 18080 25910
rect 18220 25950 18300 25960
rect 18220 25910 18240 25950
rect 18280 25910 18300 25950
rect 18220 25900 18300 25910
rect 18440 25950 18520 25960
rect 18440 25910 18460 25950
rect 18500 25910 18520 25950
rect 18440 25900 18520 25910
rect 18660 25950 18740 25960
rect 18660 25910 18680 25950
rect 18720 25910 18740 25950
rect 18660 25900 18740 25910
rect 18880 25950 18960 25960
rect 18880 25910 18900 25950
rect 18940 25910 18960 25950
rect 18880 25900 18960 25910
rect 19100 25950 19180 25960
rect 19100 25910 19120 25950
rect 19160 25910 19180 25950
rect 19100 25900 19180 25910
rect 19320 25950 19400 25960
rect 19320 25910 19340 25950
rect 19380 25910 19400 25950
rect 19320 25900 19400 25910
rect 19540 25950 19620 25960
rect 19540 25910 19560 25950
rect 19600 25910 19620 25950
rect 19540 25900 19620 25910
rect 19760 25950 19840 25960
rect 19760 25910 19780 25950
rect 19820 25910 19840 25950
rect 19760 25900 19840 25910
rect 19980 25950 20060 25960
rect 19980 25910 20000 25950
rect 20040 25910 20060 25950
rect 19980 25900 20060 25910
rect 20200 25950 20280 25960
rect 20200 25910 20220 25950
rect 20260 25910 20280 25950
rect 20200 25900 20280 25910
rect 20420 25950 20500 25960
rect 20420 25910 20440 25950
rect 20480 25910 20500 25950
rect 20420 25900 20500 25910
rect 17120 25060 17200 25070
rect 17120 25020 17140 25060
rect 17180 25020 17200 25060
rect 17120 25010 17200 25020
rect 17340 25060 17420 25070
rect 17340 25020 17360 25060
rect 17400 25020 17420 25060
rect 17340 25010 17420 25020
rect 17560 25060 17640 25070
rect 17560 25020 17580 25060
rect 17620 25020 17640 25060
rect 17560 25010 17640 25020
rect 17780 25060 17860 25070
rect 17780 25020 17800 25060
rect 17840 25020 17860 25060
rect 17780 25010 17860 25020
rect 18000 25060 18080 25070
rect 18000 25020 18020 25060
rect 18060 25020 18080 25060
rect 18000 25010 18080 25020
rect 18220 25060 18300 25070
rect 18220 25020 18240 25060
rect 18280 25020 18300 25060
rect 18220 25010 18300 25020
rect 18440 25060 18520 25070
rect 18440 25020 18460 25060
rect 18500 25020 18520 25060
rect 18440 25010 18520 25020
rect 18660 25060 18740 25070
rect 18660 25020 18680 25060
rect 18720 25020 18740 25060
rect 18660 25010 18740 25020
rect 18880 25060 18960 25070
rect 18880 25020 18900 25060
rect 18940 25020 18960 25060
rect 18880 25010 18960 25020
rect 19100 25060 19180 25070
rect 19100 25020 19120 25060
rect 19160 25020 19180 25060
rect 19100 25010 19180 25020
rect 19320 25060 19400 25070
rect 19320 25020 19340 25060
rect 19380 25020 19400 25060
rect 19320 25010 19400 25020
rect 19540 25060 19620 25070
rect 19540 25020 19560 25060
rect 19600 25020 19620 25060
rect 19540 25010 19620 25020
rect 19760 25060 19840 25070
rect 19760 25020 19780 25060
rect 19820 25020 19840 25060
rect 19760 25010 19840 25020
rect 19980 25060 20060 25070
rect 19980 25020 20000 25060
rect 20040 25020 20060 25060
rect 19980 25010 20060 25020
rect 20200 25060 20280 25070
rect 20200 25020 20220 25060
rect 20260 25020 20280 25060
rect 20200 25010 20280 25020
rect 20420 25060 20500 25070
rect 20420 25020 20440 25060
rect 20480 25020 20500 25060
rect 20420 25010 20500 25020
rect 16830 24940 16960 24950
rect 16830 24890 16890 24940
rect 16940 24890 16960 24940
rect 16830 24880 16960 24890
rect 17020 24940 17090 24960
rect 17020 24900 17040 24940
rect 17080 24900 17090 24940
rect 17020 24880 17090 24900
rect 20540 24950 20600 26020
rect 20540 24940 20670 24950
rect 20540 24890 20600 24940
rect 20650 24890 20670 24940
rect 20540 24880 20670 24890
rect 14890 24660 14900 24820
rect 14940 24660 14950 24820
rect 14890 24640 14950 24660
rect 15070 24820 15130 24840
rect 15070 24660 15080 24820
rect 15120 24660 15130 24820
rect 15070 24640 15130 24660
rect 15180 24820 15240 24840
rect 15180 24660 15190 24820
rect 15230 24660 15240 24820
rect 15180 24300 15240 24660
rect 15290 24820 15350 24840
rect 15290 24660 15300 24820
rect 15340 24660 15350 24820
rect 15290 24640 15350 24660
rect 15400 24820 15460 24840
rect 15400 24660 15410 24820
rect 15450 24660 15460 24820
rect 15400 24300 15460 24660
rect 15510 24820 15570 24840
rect 15510 24660 15520 24820
rect 15560 24660 15570 24820
rect 15510 24640 15570 24660
rect 15620 24820 15680 24840
rect 15620 24660 15630 24820
rect 15670 24660 15680 24820
rect 15620 24300 15680 24660
rect 15730 24820 15790 24840
rect 15730 24660 15740 24820
rect 15780 24660 15790 24820
rect 15730 24640 15790 24660
rect 15840 24820 15900 24840
rect 15840 24660 15850 24820
rect 15890 24660 15900 24820
rect 15840 24300 15900 24660
rect 15950 24820 16010 24840
rect 15950 24660 15960 24820
rect 16000 24660 16010 24820
rect 15950 24640 16010 24660
rect 16060 24820 16120 24840
rect 16060 24660 16070 24820
rect 16110 24660 16120 24820
rect 16060 24300 16120 24660
rect 16170 24820 16230 24840
rect 16170 24660 16180 24820
rect 16220 24660 16230 24820
rect 16170 24640 16230 24660
rect 16280 24820 16340 24840
rect 16280 24660 16290 24820
rect 16330 24660 16340 24820
rect 16280 24300 16340 24660
rect 16390 24820 16450 24840
rect 16390 24660 16400 24820
rect 16440 24660 16450 24820
rect 16390 24640 16450 24660
rect 16500 24820 16560 24840
rect 16500 24660 16510 24820
rect 16550 24660 16560 24820
rect 16500 24300 16560 24660
rect 16610 24820 16670 24840
rect 16610 24660 16620 24820
rect 16660 24660 16670 24820
rect 16610 24640 16670 24660
rect 16720 24820 16780 24840
rect 16720 24660 16730 24820
rect 16770 24660 16780 24820
rect 16720 24300 16780 24660
rect 16830 24820 16890 24880
rect 16830 24660 16840 24820
rect 16880 24660 16890 24820
rect 16830 24640 16890 24660
rect 17020 24820 17080 24840
rect 17020 24660 17030 24820
rect 17070 24660 17080 24820
rect 17020 24640 17080 24660
rect 17130 24820 17190 24840
rect 17130 24660 17140 24820
rect 17180 24660 17190 24820
rect 17130 24300 17190 24660
rect 17240 24820 17300 24840
rect 17240 24660 17250 24820
rect 17290 24660 17300 24820
rect 17240 24640 17300 24660
rect 17350 24820 17410 24840
rect 17350 24660 17360 24820
rect 17400 24660 17410 24820
rect 17350 24300 17410 24660
rect 17460 24820 17520 24840
rect 17460 24660 17470 24820
rect 17510 24660 17520 24820
rect 17460 24640 17520 24660
rect 17570 24820 17630 24840
rect 17570 24660 17580 24820
rect 17620 24660 17630 24820
rect 17570 24300 17630 24660
rect 17680 24820 17740 24840
rect 17680 24660 17690 24820
rect 17730 24660 17740 24820
rect 17680 24640 17740 24660
rect 17790 24820 17850 24840
rect 17790 24660 17800 24820
rect 17840 24660 17850 24820
rect 17790 24300 17850 24660
rect 17900 24820 17960 24840
rect 17900 24660 17910 24820
rect 17950 24660 17960 24820
rect 17900 24640 17960 24660
rect 18010 24820 18070 24840
rect 18010 24660 18020 24820
rect 18060 24660 18070 24820
rect 18010 24300 18070 24660
rect 18120 24820 18180 24840
rect 18120 24660 18130 24820
rect 18170 24660 18180 24820
rect 18120 24640 18180 24660
rect 18230 24820 18290 24840
rect 18230 24660 18240 24820
rect 18280 24660 18290 24820
rect 18230 24300 18290 24660
rect 18340 24820 18400 24840
rect 18340 24660 18350 24820
rect 18390 24660 18400 24820
rect 18340 24640 18400 24660
rect 18450 24820 18510 24840
rect 18450 24660 18460 24820
rect 18500 24660 18510 24820
rect 18450 24300 18510 24660
rect 18560 24820 18620 24840
rect 18560 24660 18570 24820
rect 18610 24660 18620 24820
rect 18560 24640 18620 24660
rect 18670 24820 18730 24840
rect 18670 24660 18680 24820
rect 18720 24660 18730 24820
rect 18670 24300 18730 24660
rect 18780 24820 18840 24840
rect 18780 24660 18790 24820
rect 18830 24660 18840 24820
rect 18780 24640 18840 24660
rect 18890 24820 18950 24840
rect 18890 24660 18900 24820
rect 18940 24660 18950 24820
rect 18890 24300 18950 24660
rect 19000 24820 19060 24840
rect 19000 24660 19010 24820
rect 19050 24660 19060 24820
rect 19000 24640 19060 24660
rect 19110 24820 19170 24840
rect 19110 24660 19120 24820
rect 19160 24660 19170 24820
rect 19110 24300 19170 24660
rect 19220 24820 19280 24840
rect 19220 24660 19230 24820
rect 19270 24660 19280 24820
rect 19220 24640 19280 24660
rect 19330 24820 19390 24840
rect 19330 24660 19340 24820
rect 19380 24660 19390 24820
rect 19330 24300 19390 24660
rect 19440 24820 19500 24840
rect 19440 24660 19450 24820
rect 19490 24660 19500 24820
rect 19440 24640 19500 24660
rect 19550 24820 19610 24840
rect 19550 24660 19560 24820
rect 19600 24660 19610 24820
rect 19550 24300 19610 24660
rect 19660 24820 19720 24840
rect 19660 24660 19670 24820
rect 19710 24660 19720 24820
rect 19660 24640 19720 24660
rect 19770 24820 19830 24840
rect 19770 24660 19780 24820
rect 19820 24660 19830 24820
rect 19770 24300 19830 24660
rect 19880 24820 19940 24840
rect 19880 24660 19890 24820
rect 19930 24660 19940 24820
rect 19880 24640 19940 24660
rect 19990 24820 20050 24840
rect 19990 24660 20000 24820
rect 20040 24660 20050 24820
rect 19990 24300 20050 24660
rect 20100 24820 20160 24840
rect 20100 24660 20110 24820
rect 20150 24660 20160 24820
rect 20100 24640 20160 24660
rect 20210 24820 20270 24840
rect 20210 24660 20220 24820
rect 20260 24660 20270 24820
rect 20210 24300 20270 24660
rect 20320 24820 20380 24840
rect 20320 24660 20330 24820
rect 20370 24660 20380 24820
rect 20320 24640 20380 24660
rect 20430 24820 20490 24840
rect 20430 24660 20440 24820
rect 20480 24660 20490 24820
rect 20430 24300 20490 24660
rect 20540 24820 20600 24880
rect 20540 24660 20550 24820
rect 20590 24660 20600 24820
rect 20540 24640 20600 24660
rect 7280 24290 20620 24300
rect 7280 24250 7320 24290
rect 7360 24250 7400 24290
rect 7440 24250 7480 24290
rect 7520 24250 7560 24290
rect 7600 24250 7640 24290
rect 7680 24250 7720 24290
rect 7760 24250 7800 24290
rect 7840 24250 7890 24290
rect 7930 24250 7970 24290
rect 8010 24250 8050 24290
rect 8090 24250 8130 24290
rect 8170 24250 8210 24290
rect 8250 24250 8290 24290
rect 8330 24250 8400 24290
rect 8440 24250 8520 24290
rect 8560 24250 8600 24290
rect 8640 24250 8680 24290
rect 8720 24250 8760 24290
rect 8800 24250 8840 24290
rect 8880 24250 8920 24290
rect 8960 24250 9000 24290
rect 9040 24250 9080 24290
rect 9120 24250 9160 24290
rect 9200 24250 9270 24290
rect 9310 24250 9350 24290
rect 9390 24250 9430 24290
rect 9470 24250 9510 24290
rect 9550 24250 9590 24290
rect 9630 24250 9670 24290
rect 9710 24250 9750 24290
rect 9790 24250 9830 24290
rect 9870 24250 9910 24290
rect 9950 24250 9990 24290
rect 10030 24250 10070 24290
rect 10110 24250 10150 24290
rect 10190 24250 10230 24290
rect 10270 24250 10310 24290
rect 10350 24250 10390 24290
rect 10430 24250 10470 24290
rect 10510 24250 10550 24290
rect 10590 24250 10630 24290
rect 10670 24250 10710 24290
rect 10750 24250 10790 24290
rect 10830 24250 10870 24290
rect 10910 24250 10950 24290
rect 10990 24250 11030 24290
rect 11070 24250 11110 24290
rect 11150 24250 11190 24290
rect 11230 24250 11270 24290
rect 11310 24250 11350 24290
rect 11390 24250 11430 24290
rect 11470 24250 11510 24290
rect 11550 24250 11590 24290
rect 11630 24250 11670 24290
rect 11710 24250 11750 24290
rect 11790 24250 11830 24290
rect 11870 24250 11910 24290
rect 11950 24250 11990 24290
rect 12030 24250 12070 24290
rect 12110 24250 12150 24290
rect 12190 24250 12230 24290
rect 12270 24250 12310 24290
rect 12350 24250 12390 24290
rect 12430 24250 12470 24290
rect 12510 24250 12550 24290
rect 12590 24250 12630 24290
rect 12670 24250 12710 24290
rect 12750 24250 12790 24290
rect 12830 24250 12870 24290
rect 12910 24250 12950 24290
rect 12990 24250 13030 24290
rect 13070 24250 13110 24290
rect 13150 24250 13190 24290
rect 13230 24250 13270 24290
rect 13310 24250 13350 24290
rect 13390 24250 13430 24290
rect 13470 24250 13510 24290
rect 13550 24250 13590 24290
rect 13630 24250 13670 24290
rect 13710 24250 13750 24290
rect 13790 24250 13830 24290
rect 13870 24250 13910 24290
rect 13950 24250 13990 24290
rect 14030 24250 14070 24290
rect 14110 24250 14150 24290
rect 14190 24250 14230 24290
rect 14270 24250 14310 24290
rect 14350 24250 14390 24290
rect 14430 24250 14470 24290
rect 14510 24250 14550 24290
rect 14590 24250 14630 24290
rect 14670 24250 14710 24290
rect 14750 24250 14790 24290
rect 14830 24250 14870 24290
rect 14910 24250 14950 24290
rect 14990 24250 15030 24290
rect 15070 24250 15110 24290
rect 15150 24250 15190 24290
rect 15230 24250 15270 24290
rect 15310 24250 15350 24290
rect 15390 24250 15430 24290
rect 15470 24250 15510 24290
rect 15550 24250 15590 24290
rect 15630 24250 15670 24290
rect 15710 24250 15750 24290
rect 15790 24250 15830 24290
rect 15870 24250 15910 24290
rect 15950 24250 15990 24290
rect 16030 24250 16070 24290
rect 16110 24250 16150 24290
rect 16190 24250 16230 24290
rect 16270 24250 16310 24290
rect 16350 24250 16390 24290
rect 16430 24250 16470 24290
rect 16510 24250 16550 24290
rect 16590 24250 16630 24290
rect 16670 24250 16710 24290
rect 16750 24250 16790 24290
rect 16830 24250 16870 24290
rect 16910 24250 16950 24290
rect 16990 24250 17030 24290
rect 17070 24250 17110 24290
rect 17150 24250 17190 24290
rect 17230 24250 17270 24290
rect 17310 24250 17350 24290
rect 17390 24250 17430 24290
rect 17470 24250 17510 24290
rect 17550 24250 17590 24290
rect 17630 24250 17670 24290
rect 17710 24250 17750 24290
rect 17790 24250 17830 24290
rect 17870 24250 17910 24290
rect 17950 24250 17990 24290
rect 18030 24250 18070 24290
rect 18110 24250 18150 24290
rect 18190 24250 18230 24290
rect 18270 24250 18310 24290
rect 18350 24250 18390 24290
rect 18430 24250 18470 24290
rect 18510 24250 18550 24290
rect 18590 24250 18630 24290
rect 18670 24250 18710 24290
rect 18750 24250 18790 24290
rect 18830 24250 18870 24290
rect 18910 24250 18950 24290
rect 18990 24250 19030 24290
rect 19070 24250 19110 24290
rect 19150 24250 19190 24290
rect 19230 24250 19270 24290
rect 19310 24250 19350 24290
rect 19390 24250 19430 24290
rect 19470 24250 19510 24290
rect 19550 24250 19590 24290
rect 19630 24250 19670 24290
rect 19710 24250 19750 24290
rect 19790 24250 19830 24290
rect 19870 24250 19910 24290
rect 19950 24250 19990 24290
rect 20030 24250 20070 24290
rect 20110 24250 20150 24290
rect 20190 24250 20230 24290
rect 20270 24250 20310 24290
rect 20350 24250 20390 24290
rect 20430 24250 20470 24290
rect 20510 24250 20550 24290
rect 20590 24250 20620 24290
rect 7280 24240 20620 24250
rect 7280 23320 20620 23330
rect 7280 23280 7310 23320
rect 7350 23280 7390 23320
rect 7430 23280 7470 23320
rect 7510 23280 7550 23320
rect 7590 23280 7630 23320
rect 7670 23280 7710 23320
rect 7750 23280 7790 23320
rect 7830 23280 7870 23320
rect 7910 23280 7950 23320
rect 7990 23280 8030 23320
rect 8070 23280 8110 23320
rect 8150 23280 8190 23320
rect 8230 23280 8270 23320
rect 8310 23280 8350 23320
rect 8390 23280 8430 23320
rect 8470 23280 8520 23320
rect 8560 23280 8600 23320
rect 8640 23280 8680 23320
rect 8720 23280 8760 23320
rect 8800 23280 8840 23320
rect 8880 23280 8920 23320
rect 8960 23280 9000 23320
rect 9040 23280 9080 23320
rect 9120 23280 9160 23320
rect 9200 23280 9270 23320
rect 9310 23280 9350 23320
rect 9390 23280 9430 23320
rect 9470 23280 9510 23320
rect 9550 23280 9590 23320
rect 9630 23280 9670 23320
rect 9710 23280 9750 23320
rect 9790 23280 9830 23320
rect 9870 23280 9910 23320
rect 9950 23280 9990 23320
rect 10030 23280 10070 23320
rect 10110 23280 10150 23320
rect 10190 23280 10230 23320
rect 10270 23280 10310 23320
rect 10350 23280 10390 23320
rect 10430 23280 10470 23320
rect 10510 23280 10550 23320
rect 10590 23280 10630 23320
rect 10670 23280 10710 23320
rect 10750 23280 10790 23320
rect 10830 23280 10870 23320
rect 10910 23280 10950 23320
rect 10990 23280 11030 23320
rect 11070 23280 11110 23320
rect 11150 23280 11190 23320
rect 11230 23280 11270 23320
rect 11310 23280 11350 23320
rect 11390 23280 11430 23320
rect 11470 23280 11510 23320
rect 11550 23280 11590 23320
rect 11630 23280 11670 23320
rect 11710 23280 11750 23320
rect 11790 23280 11830 23320
rect 11870 23280 11910 23320
rect 11950 23280 11990 23320
rect 12030 23280 12070 23320
rect 12110 23280 12150 23320
rect 12190 23280 12230 23320
rect 12270 23280 12310 23320
rect 12350 23280 12390 23320
rect 12430 23280 12470 23320
rect 12510 23280 12550 23320
rect 12590 23280 12630 23320
rect 12670 23280 12710 23320
rect 12750 23280 12790 23320
rect 12830 23280 12870 23320
rect 12910 23280 12950 23320
rect 12990 23280 13030 23320
rect 13070 23280 13110 23320
rect 13150 23280 13190 23320
rect 13230 23280 13270 23320
rect 13310 23280 13350 23320
rect 13390 23280 13430 23320
rect 13470 23280 13510 23320
rect 13550 23280 13590 23320
rect 13630 23280 13670 23320
rect 13710 23280 13750 23320
rect 13790 23280 13830 23320
rect 13870 23280 13910 23320
rect 13950 23280 13990 23320
rect 14030 23280 14070 23320
rect 14110 23280 14150 23320
rect 14190 23280 14230 23320
rect 14270 23280 14310 23320
rect 14350 23280 14390 23320
rect 14430 23280 14470 23320
rect 14510 23280 14550 23320
rect 14590 23280 14630 23320
rect 14670 23280 14710 23320
rect 14750 23280 14790 23320
rect 14830 23280 14870 23320
rect 14910 23280 14950 23320
rect 14990 23280 15030 23320
rect 15070 23280 15110 23320
rect 15150 23280 15190 23320
rect 15230 23280 15270 23320
rect 15310 23280 15350 23320
rect 15390 23280 15430 23320
rect 15470 23280 15510 23320
rect 15550 23280 15590 23320
rect 15630 23280 15670 23320
rect 15710 23280 15750 23320
rect 15790 23280 15830 23320
rect 15870 23280 15910 23320
rect 15950 23280 15990 23320
rect 16030 23280 16070 23320
rect 16110 23280 16150 23320
rect 16190 23280 16230 23320
rect 16270 23280 16310 23320
rect 16350 23280 16390 23320
rect 16430 23280 16470 23320
rect 16510 23280 16550 23320
rect 16590 23280 16630 23320
rect 16670 23280 16710 23320
rect 16750 23280 16790 23320
rect 16830 23280 16870 23320
rect 16910 23280 16950 23320
rect 16990 23280 17030 23320
rect 17070 23280 17110 23320
rect 17150 23280 17190 23320
rect 17230 23280 17270 23320
rect 17310 23280 17350 23320
rect 17390 23280 17430 23320
rect 17470 23280 17510 23320
rect 17550 23280 17590 23320
rect 17630 23280 17670 23320
rect 17710 23280 17750 23320
rect 17790 23280 17830 23320
rect 17870 23280 17910 23320
rect 17950 23280 17990 23320
rect 18030 23280 18070 23320
rect 18110 23280 18150 23320
rect 18190 23280 18230 23320
rect 18270 23280 18310 23320
rect 18350 23280 18390 23320
rect 18430 23280 18470 23320
rect 18510 23280 18550 23320
rect 18590 23280 18630 23320
rect 18670 23280 18710 23320
rect 18750 23280 18790 23320
rect 18830 23280 18870 23320
rect 18910 23280 18950 23320
rect 18990 23280 19030 23320
rect 19070 23280 19110 23320
rect 19150 23280 19190 23320
rect 19230 23280 19270 23320
rect 19310 23280 19350 23320
rect 19390 23280 19430 23320
rect 19470 23280 19510 23320
rect 19550 23280 19590 23320
rect 19630 23280 19670 23320
rect 19710 23280 19750 23320
rect 19790 23280 19830 23320
rect 19870 23280 19910 23320
rect 19950 23280 19990 23320
rect 20030 23280 20070 23320
rect 20110 23280 20150 23320
rect 20190 23280 20230 23320
rect 20270 23280 20310 23320
rect 20350 23280 20390 23320
rect 20430 23280 20470 23320
rect 20510 23280 20550 23320
rect 20590 23280 20620 23320
rect 7280 23270 20620 23280
rect 7470 23190 7530 23270
rect 7470 22830 7480 23190
rect 7520 22830 7530 23190
rect 7470 22810 7530 22830
rect 7730 23190 7790 23210
rect 7730 22830 7740 23190
rect 7780 22830 7790 23190
rect 7960 23190 8020 23270
rect 7960 23030 7970 23190
rect 8010 23030 8020 23190
rect 7960 23010 8020 23030
rect 8070 23190 8130 23210
rect 8070 23030 8080 23190
rect 8120 23030 8130 23190
rect 7630 22770 7690 22790
rect 7630 22730 7640 22770
rect 7680 22730 7690 22770
rect 7630 22710 7690 22730
rect 7370 22680 7430 22700
rect 7370 22640 7380 22680
rect 7420 22640 7430 22680
rect 7730 22680 7790 22830
rect 8070 22680 8130 23030
rect 8180 23190 8240 23270
rect 8180 23030 8190 23190
rect 8230 23030 8240 23190
rect 8180 23010 8240 23030
rect 8480 23190 8540 23270
rect 8480 22830 8490 23190
rect 8530 22830 8540 23190
rect 8480 22810 8540 22830
rect 8610 23190 8670 23210
rect 8610 22830 8620 23190
rect 8660 22830 8670 23190
rect 8610 22810 8670 22830
rect 8740 23190 8800 23210
rect 8740 22830 8750 23190
rect 8790 22830 8800 23190
rect 8630 22750 8700 22770
rect 8630 22710 8650 22750
rect 8690 22710 8700 22750
rect 8630 22690 8700 22710
rect 8740 22690 8800 22830
rect 8860 22920 8920 23270
rect 9220 23190 9280 23270
rect 9220 23030 9230 23190
rect 9270 23030 9280 23190
rect 9220 23010 9280 23030
rect 9330 23190 9390 23210
rect 9330 23030 9340 23190
rect 9380 23030 9390 23190
rect 8860 22760 8870 22920
rect 8910 22760 8920 22920
rect 8860 22740 8920 22760
rect 8970 22920 9030 22940
rect 8970 22760 8980 22920
rect 9020 22760 9030 22920
rect 9080 22910 9170 22930
rect 9080 22860 9100 22910
rect 9150 22860 9170 22910
rect 9080 22840 9170 22860
rect 8970 22690 9030 22760
rect 9090 22690 9160 22840
rect 9330 22770 9390 23030
rect 9440 23190 9500 23270
rect 9440 23030 9450 23190
rect 9490 23030 9500 23190
rect 9440 23010 9500 23030
rect 9670 23190 9730 23270
rect 9670 22830 9680 23190
rect 9720 22830 9730 23190
rect 9670 22810 9730 22830
rect 9930 23190 9990 23210
rect 9930 22830 9940 23190
rect 9980 22830 9990 23190
rect 10160 23190 10220 23270
rect 10160 23030 10170 23190
rect 10210 23030 10220 23190
rect 10160 23010 10220 23030
rect 10270 23190 10330 23210
rect 10270 23030 10280 23190
rect 10320 23030 10330 23190
rect 9830 22770 9890 22790
rect 9330 22730 9840 22770
rect 9880 22730 9890 22770
rect 7730 22670 8030 22680
rect 7370 22620 7430 22640
rect 7600 22630 7880 22670
rect 7920 22630 7960 22670
rect 8000 22630 8030 22670
rect 7600 22620 8030 22630
rect 8070 22670 8320 22680
rect 8070 22630 8260 22670
rect 8300 22630 8320 22670
rect 8070 22620 8320 22630
rect 8480 22670 8550 22690
rect 8480 22630 8500 22670
rect 8540 22630 8550 22670
rect 8740 22670 8930 22690
rect 8740 22650 8800 22670
rect 7460 22560 7540 22570
rect 7460 22520 7480 22560
rect 7520 22520 7540 22560
rect 7460 22510 7540 22520
rect 7460 21700 7540 21710
rect 7460 21660 7480 21700
rect 7520 21660 7540 21700
rect 7460 21650 7540 21660
rect 7470 21560 7530 21580
rect 7470 21100 7480 21560
rect 7520 21100 7530 21560
rect 7470 21010 7530 21100
rect 7600 21560 7660 22620
rect 7720 22560 7800 22570
rect 7720 22520 7740 22560
rect 7780 22520 7800 22560
rect 7720 22510 7800 22520
rect 7720 21680 7800 21690
rect 7720 21640 7740 21680
rect 7780 21640 7800 21680
rect 7720 21630 7800 21640
rect 7600 21100 7610 21560
rect 7650 21100 7660 21560
rect 7600 21080 7660 21100
rect 7730 21560 7790 21580
rect 7730 21100 7740 21560
rect 7780 21100 7790 21560
rect 7730 21010 7790 21100
rect 7960 21560 8020 21580
rect 7960 21100 7970 21560
rect 8010 21100 8020 21560
rect 7960 21010 8020 21100
rect 8070 21560 8130 22620
rect 8480 22610 8550 22630
rect 8610 22630 8800 22650
rect 8840 22630 8880 22670
rect 8920 22630 8930 22670
rect 8610 22610 8930 22630
rect 8970 22670 9160 22690
rect 8970 22630 9000 22670
rect 9040 22630 9160 22670
rect 8970 22610 9160 22630
rect 9200 22700 9290 22720
rect 9200 22640 9220 22700
rect 9280 22640 9290 22700
rect 9200 22620 9290 22640
rect 8070 21100 8080 21560
rect 8120 21100 8130 21560
rect 8070 21080 8130 21100
rect 8180 21560 8240 21580
rect 8180 21100 8190 21560
rect 8230 21100 8240 21560
rect 8180 21010 8240 21100
rect 8480 21550 8540 21570
rect 8480 21090 8490 21550
rect 8530 21090 8540 21550
rect 8480 21010 8540 21090
rect 8610 21550 8670 22610
rect 8610 21090 8620 21550
rect 8660 21090 8670 21550
rect 8610 21070 8670 21090
rect 8740 21550 8800 21570
rect 8740 21090 8750 21550
rect 8790 21090 8800 21550
rect 8740 21010 8800 21090
rect 8860 21550 8920 21570
rect 8860 21090 8870 21550
rect 8910 21090 8920 21550
rect 8860 21010 8920 21090
rect 8970 21550 9030 22610
rect 8970 21090 8980 21550
rect 9020 21090 9030 21550
rect 8970 21070 9030 21090
rect 9220 21550 9280 21570
rect 9220 21090 9230 21550
rect 9270 21090 9280 21550
rect 9220 21010 9280 21090
rect 9330 21550 9390 22730
rect 9830 22710 9890 22730
rect 9570 22670 9630 22690
rect 9930 22670 9990 22830
rect 10270 22670 10330 23030
rect 10380 23190 10440 23270
rect 10380 23030 10390 23190
rect 10430 23030 10440 23190
rect 10380 23010 10440 23030
rect 10660 23190 10720 23270
rect 10660 22830 10670 23190
rect 10710 22830 10720 23190
rect 10660 22810 10720 22830
rect 10920 23190 10980 23210
rect 10920 22830 10930 23190
rect 10970 22830 10980 23190
rect 11150 23190 11210 23270
rect 11150 23030 11160 23190
rect 11200 23030 11210 23190
rect 11150 23010 11210 23030
rect 11260 23190 11320 23210
rect 11260 23030 11270 23190
rect 11310 23030 11320 23190
rect 10820 22770 10880 22790
rect 10820 22730 10830 22770
rect 10870 22730 10880 22770
rect 10820 22710 10880 22730
rect 10560 22670 10620 22690
rect 10920 22670 10980 22830
rect 11260 22670 11320 23030
rect 11370 23190 11430 23270
rect 11370 23030 11380 23190
rect 11420 23030 11430 23190
rect 11370 23010 11430 23030
rect 11660 23190 11720 23270
rect 11660 22830 11670 23190
rect 11710 22830 11720 23190
rect 11660 22810 11720 22830
rect 11920 23190 11980 23210
rect 11920 22830 11930 23190
rect 11970 22830 11980 23190
rect 12150 23190 12210 23270
rect 12150 23030 12160 23190
rect 12200 23030 12210 23190
rect 12150 23010 12210 23030
rect 12260 23190 12320 23210
rect 12260 23030 12270 23190
rect 12310 23030 12320 23190
rect 11820 22770 11880 22790
rect 11820 22730 11830 22770
rect 11870 22730 11880 22770
rect 11820 22710 11880 22730
rect 11560 22670 11620 22690
rect 11920 22670 11980 22830
rect 12260 22670 12320 23030
rect 12370 23190 12430 23270
rect 12370 23030 12380 23190
rect 12420 23030 12430 23190
rect 12370 23010 12430 23030
rect 12530 23190 12590 23270
rect 12530 23030 12540 23190
rect 12580 23030 12590 23190
rect 12530 23010 12590 23030
rect 12640 23190 12700 23210
rect 12640 23030 12650 23190
rect 12690 23030 12700 23190
rect 12640 22690 12700 23030
rect 12750 23190 12810 23270
rect 12750 23030 12760 23190
rect 12800 23030 12810 23190
rect 12750 23010 12810 23030
rect 12880 22910 12940 23270
rect 12880 22750 12890 22910
rect 12930 22750 12940 22910
rect 12880 22730 12940 22750
rect 12990 22910 13050 22930
rect 12990 22750 13000 22910
rect 13040 22750 13050 22910
rect 12640 22670 12950 22690
rect 9570 22630 9580 22670
rect 9620 22630 9630 22670
rect 9570 22610 9630 22630
rect 9800 22660 10230 22670
rect 9800 22620 10080 22660
rect 10120 22620 10160 22660
rect 10200 22620 10230 22660
rect 9800 22610 10230 22620
rect 10270 22660 10510 22670
rect 10270 22620 10460 22660
rect 10500 22620 10510 22660
rect 10270 22610 10510 22620
rect 10560 22630 10570 22670
rect 10610 22630 10620 22670
rect 10560 22610 10620 22630
rect 10790 22660 11220 22670
rect 10790 22620 11070 22660
rect 11110 22620 11150 22660
rect 11190 22620 11220 22660
rect 10790 22610 11220 22620
rect 11260 22660 11500 22670
rect 11260 22620 11450 22660
rect 11490 22620 11500 22660
rect 11260 22610 11500 22620
rect 11560 22630 11570 22670
rect 11610 22630 11620 22670
rect 11560 22610 11620 22630
rect 11790 22660 12220 22670
rect 11790 22620 12070 22660
rect 12110 22620 12150 22660
rect 12190 22620 12220 22660
rect 11790 22610 12220 22620
rect 12260 22660 12600 22670
rect 12260 22620 12450 22660
rect 12490 22620 12530 22660
rect 12570 22620 12600 22660
rect 12260 22610 12600 22620
rect 12640 22630 12820 22670
rect 12860 22630 12900 22670
rect 12940 22630 12950 22670
rect 12640 22610 12950 22630
rect 12990 22670 13050 22750
rect 13110 22910 13170 22930
rect 13110 22750 13120 22910
rect 13160 22750 13170 22910
rect 13110 22730 13170 22750
rect 13220 22910 13280 23270
rect 13220 22750 13230 22910
rect 13270 22750 13280 22910
rect 13220 22730 13280 22750
rect 13330 22910 13390 22930
rect 13330 22750 13340 22910
rect 13380 22750 13390 22910
rect 12990 22630 13000 22670
rect 13040 22630 13050 22670
rect 9660 22550 9740 22560
rect 9660 22510 9680 22550
rect 9720 22510 9740 22550
rect 9660 22500 9740 22510
rect 9660 21670 9740 21680
rect 9660 21630 9680 21670
rect 9720 21630 9740 21670
rect 9660 21620 9740 21630
rect 9330 21090 9340 21550
rect 9380 21090 9390 21550
rect 9330 21070 9390 21090
rect 9440 21550 9500 21570
rect 9440 21090 9450 21550
rect 9490 21090 9500 21550
rect 9440 21010 9500 21090
rect 9670 21550 9730 21570
rect 9670 21090 9680 21550
rect 9720 21090 9730 21550
rect 9670 21010 9730 21090
rect 9800 21550 9860 22610
rect 9920 22550 10000 22560
rect 9920 22510 9940 22550
rect 9980 22510 10000 22550
rect 9920 22500 10000 22510
rect 9920 21670 10000 21680
rect 9920 21630 9940 21670
rect 9980 21630 10000 21670
rect 9920 21620 10000 21630
rect 9800 21090 9810 21550
rect 9850 21090 9860 21550
rect 9800 21070 9860 21090
rect 9930 21550 9990 21570
rect 9930 21090 9940 21550
rect 9980 21090 9990 21550
rect 9930 21010 9990 21090
rect 10160 21550 10220 21570
rect 10160 21090 10170 21550
rect 10210 21090 10220 21550
rect 10160 21010 10220 21090
rect 10270 21550 10330 22610
rect 10650 22550 10730 22560
rect 10650 22510 10670 22550
rect 10710 22510 10730 22550
rect 10650 22500 10730 22510
rect 10650 21670 10730 21680
rect 10650 21630 10670 21670
rect 10710 21630 10730 21670
rect 10650 21620 10730 21630
rect 10270 21090 10280 21550
rect 10320 21090 10330 21550
rect 10270 21070 10330 21090
rect 10380 21550 10440 21570
rect 10380 21090 10390 21550
rect 10430 21090 10440 21550
rect 10380 21010 10440 21090
rect 10660 21550 10720 21570
rect 10660 21090 10670 21550
rect 10710 21090 10720 21550
rect 10660 21010 10720 21090
rect 10790 21550 10850 22610
rect 10910 22550 10990 22560
rect 10910 22510 10930 22550
rect 10970 22510 10990 22550
rect 10910 22500 10990 22510
rect 10910 21670 10990 21680
rect 10910 21630 10930 21670
rect 10970 21630 10990 21670
rect 10910 21620 10990 21630
rect 10790 21090 10800 21550
rect 10840 21090 10850 21550
rect 10790 21070 10850 21090
rect 10920 21550 10980 21570
rect 10920 21090 10930 21550
rect 10970 21090 10980 21550
rect 10920 21010 10980 21090
rect 11150 21550 11210 21570
rect 11150 21090 11160 21550
rect 11200 21090 11210 21550
rect 11150 21010 11210 21090
rect 11260 21550 11320 22610
rect 11650 22550 11730 22560
rect 11650 22510 11670 22550
rect 11710 22510 11730 22550
rect 11650 22500 11730 22510
rect 11650 21670 11730 21680
rect 11650 21630 11670 21670
rect 11710 21630 11730 21670
rect 11650 21620 11730 21630
rect 11260 21090 11270 21550
rect 11310 21090 11320 21550
rect 11260 21070 11320 21090
rect 11370 21550 11430 21570
rect 11370 21090 11380 21550
rect 11420 21090 11430 21550
rect 11370 21010 11430 21090
rect 11660 21550 11720 21570
rect 11660 21090 11670 21550
rect 11710 21090 11720 21550
rect 11660 21010 11720 21090
rect 11790 21550 11850 22610
rect 11910 22550 11990 22560
rect 11910 22510 11930 22550
rect 11970 22510 11990 22550
rect 11910 22500 11990 22510
rect 11910 21670 11990 21680
rect 11910 21630 11930 21670
rect 11970 21630 11990 21670
rect 11910 21620 11990 21630
rect 11790 21090 11800 21550
rect 11840 21090 11850 21550
rect 11790 21070 11850 21090
rect 11920 21550 11980 21570
rect 11920 21090 11930 21550
rect 11970 21090 11980 21550
rect 11920 21010 11980 21090
rect 12150 21550 12210 21570
rect 12150 21090 12160 21550
rect 12200 21090 12210 21550
rect 12150 21010 12210 21090
rect 12260 21550 12320 22610
rect 12260 21090 12270 21550
rect 12310 21090 12320 21550
rect 12260 21070 12320 21090
rect 12370 21550 12430 21570
rect 12370 21090 12380 21550
rect 12420 21090 12430 21550
rect 12370 21010 12430 21090
rect 12530 21550 12590 21570
rect 12530 21090 12540 21550
rect 12580 21090 12590 21550
rect 12530 21010 12590 21090
rect 12640 21550 12700 22610
rect 12640 21090 12650 21550
rect 12690 21090 12700 21550
rect 12640 21070 12700 21090
rect 12750 21550 12810 21570
rect 12750 21090 12760 21550
rect 12800 21090 12810 21550
rect 12750 21010 12810 21090
rect 12880 21550 12940 21570
rect 12880 21090 12890 21550
rect 12930 21090 12940 21550
rect 12880 21010 12940 21090
rect 12990 21550 13050 22630
rect 13120 22670 13180 22690
rect 13120 22630 13130 22670
rect 13170 22630 13180 22670
rect 13120 22610 13180 22630
rect 13330 22670 13390 22750
rect 13450 22910 13510 22930
rect 13450 22750 13460 22910
rect 13500 22750 13510 22910
rect 13450 22730 13510 22750
rect 13560 22910 13620 23270
rect 13560 22750 13570 22910
rect 13610 22750 13620 22910
rect 13560 22730 13620 22750
rect 13670 22910 13730 22930
rect 13670 22750 13680 22910
rect 13720 22750 13730 22910
rect 13670 22730 13730 22750
rect 13780 22910 13840 23270
rect 13780 22750 13790 22910
rect 13830 22750 13840 22910
rect 13780 22730 13840 22750
rect 13890 22910 13950 22930
rect 13890 22750 13900 22910
rect 13940 22750 13950 22910
rect 13330 22630 13340 22670
rect 13380 22630 13390 22670
rect 13210 22570 13290 22580
rect 13210 22530 13230 22570
rect 13270 22530 13290 22570
rect 13210 22520 13290 22530
rect 13210 21680 13290 21690
rect 13210 21640 13230 21680
rect 13270 21640 13290 21680
rect 13210 21630 13290 21640
rect 12990 21090 13000 21550
rect 13040 21090 13050 21550
rect 12990 21070 13050 21090
rect 13110 21550 13170 21570
rect 13110 21090 13120 21550
rect 13160 21090 13170 21550
rect 13110 21070 13170 21090
rect 13220 21550 13280 21570
rect 13220 21090 13230 21550
rect 13270 21090 13280 21550
rect 13220 21010 13280 21090
rect 13330 21550 13390 22630
rect 13460 22670 13520 22690
rect 13460 22630 13470 22670
rect 13510 22630 13520 22670
rect 13460 22610 13520 22630
rect 13890 22670 13950 22750
rect 14010 22910 14070 22930
rect 14010 22750 14020 22910
rect 14060 22750 14070 22910
rect 14010 22730 14070 22750
rect 14120 22910 14180 23270
rect 14120 22750 14130 22910
rect 14170 22750 14180 22910
rect 14120 22730 14180 22750
rect 14230 22910 14290 22930
rect 14230 22750 14240 22910
rect 14280 22750 14290 22910
rect 14230 22730 14290 22750
rect 14340 22910 14400 23270
rect 14340 22750 14350 22910
rect 14390 22750 14400 22910
rect 14340 22730 14400 22750
rect 14450 22910 14510 22930
rect 14450 22750 14460 22910
rect 14500 22750 14510 22910
rect 14450 22730 14510 22750
rect 14560 22910 14620 23270
rect 14560 22750 14570 22910
rect 14610 22750 14620 22910
rect 14560 22730 14620 22750
rect 14670 22910 14730 22930
rect 14670 22750 14680 22910
rect 14720 22750 14730 22910
rect 14670 22730 14730 22750
rect 14780 22910 14840 23270
rect 14780 22750 14790 22910
rect 14830 22750 14840 22910
rect 14780 22730 14840 22750
rect 14890 22910 14950 22930
rect 14890 22750 14900 22910
rect 14940 22750 14950 22910
rect 13890 22630 13900 22670
rect 13940 22630 13950 22670
rect 13550 22570 13630 22580
rect 13550 22530 13570 22570
rect 13610 22530 13630 22570
rect 13550 22520 13630 22530
rect 13770 22570 13850 22580
rect 13770 22530 13790 22570
rect 13830 22530 13850 22570
rect 13770 22520 13850 22530
rect 13550 21680 13630 21690
rect 13550 21640 13570 21680
rect 13610 21640 13630 21680
rect 13550 21630 13630 21640
rect 13770 21680 13850 21690
rect 13770 21640 13790 21680
rect 13830 21640 13850 21680
rect 13770 21630 13850 21640
rect 13330 21090 13340 21550
rect 13380 21090 13390 21550
rect 13330 21070 13390 21090
rect 13450 21550 13510 21570
rect 13450 21090 13460 21550
rect 13500 21090 13510 21550
rect 13450 21070 13510 21090
rect 13560 21550 13620 21570
rect 13560 21090 13570 21550
rect 13610 21090 13620 21550
rect 13560 21010 13620 21090
rect 13670 21550 13730 21570
rect 13670 21090 13680 21550
rect 13720 21090 13730 21550
rect 13670 21070 13730 21090
rect 13780 21550 13840 21570
rect 13780 21090 13790 21550
rect 13830 21090 13840 21550
rect 13780 21010 13840 21090
rect 13890 21550 13950 22630
rect 14020 22670 14080 22690
rect 14020 22630 14030 22670
rect 14070 22630 14080 22670
rect 14020 22610 14080 22630
rect 14890 22670 14950 22750
rect 15070 22910 15130 22930
rect 15070 22750 15080 22910
rect 15120 22750 15130 22910
rect 15070 22730 15130 22750
rect 15180 22910 15240 23270
rect 15180 22750 15190 22910
rect 15230 22750 15240 22910
rect 15180 22730 15240 22750
rect 15290 22910 15350 22930
rect 15290 22750 15300 22910
rect 15340 22750 15350 22910
rect 15290 22730 15350 22750
rect 15400 22910 15460 23270
rect 15400 22750 15410 22910
rect 15450 22750 15460 22910
rect 15400 22730 15460 22750
rect 15510 22910 15570 22930
rect 15510 22750 15520 22910
rect 15560 22750 15570 22910
rect 15510 22730 15570 22750
rect 15620 22910 15680 23270
rect 15620 22750 15630 22910
rect 15670 22750 15680 22910
rect 15620 22730 15680 22750
rect 15730 22910 15790 22930
rect 15730 22750 15740 22910
rect 15780 22750 15790 22910
rect 15730 22730 15790 22750
rect 15840 22910 15900 23270
rect 15840 22750 15850 22910
rect 15890 22750 15900 22910
rect 15840 22730 15900 22750
rect 15950 22910 16010 22930
rect 15950 22750 15960 22910
rect 16000 22750 16010 22910
rect 15950 22730 16010 22750
rect 16060 22910 16120 23270
rect 16060 22750 16070 22910
rect 16110 22750 16120 22910
rect 16060 22730 16120 22750
rect 16170 22910 16230 22930
rect 16170 22750 16180 22910
rect 16220 22750 16230 22910
rect 16170 22730 16230 22750
rect 16280 22910 16340 23270
rect 16280 22750 16290 22910
rect 16330 22750 16340 22910
rect 16280 22730 16340 22750
rect 16390 22910 16450 22930
rect 16390 22750 16400 22910
rect 16440 22750 16450 22910
rect 16390 22730 16450 22750
rect 16500 22910 16560 23270
rect 16500 22750 16510 22910
rect 16550 22750 16560 22910
rect 16500 22730 16560 22750
rect 16610 22910 16670 22930
rect 16610 22750 16620 22910
rect 16660 22750 16670 22910
rect 16610 22730 16670 22750
rect 16720 22910 16780 23270
rect 16720 22750 16730 22910
rect 16770 22750 16780 22910
rect 16720 22730 16780 22750
rect 16830 22910 16890 22930
rect 16830 22750 16840 22910
rect 16880 22750 16890 22910
rect 16830 22690 16890 22750
rect 17020 22910 17080 22930
rect 17020 22750 17030 22910
rect 17070 22750 17080 22910
rect 17020 22730 17080 22750
rect 17130 22910 17190 23270
rect 17130 22750 17140 22910
rect 17180 22750 17190 22910
rect 17130 22730 17190 22750
rect 17240 22910 17300 22930
rect 17240 22750 17250 22910
rect 17290 22750 17300 22910
rect 17240 22730 17300 22750
rect 17350 22910 17410 23270
rect 17350 22750 17360 22910
rect 17400 22750 17410 22910
rect 17350 22730 17410 22750
rect 17460 22910 17520 22930
rect 17460 22750 17470 22910
rect 17510 22750 17520 22910
rect 17460 22730 17520 22750
rect 17570 22910 17630 23270
rect 17570 22750 17580 22910
rect 17620 22750 17630 22910
rect 17570 22730 17630 22750
rect 17680 22910 17740 22930
rect 17680 22750 17690 22910
rect 17730 22750 17740 22910
rect 17680 22730 17740 22750
rect 17790 22910 17850 23270
rect 17790 22750 17800 22910
rect 17840 22750 17850 22910
rect 17790 22730 17850 22750
rect 17900 22910 17960 22930
rect 17900 22750 17910 22910
rect 17950 22750 17960 22910
rect 17900 22730 17960 22750
rect 18010 22910 18070 23270
rect 18010 22750 18020 22910
rect 18060 22750 18070 22910
rect 18010 22730 18070 22750
rect 18120 22910 18180 22930
rect 18120 22750 18130 22910
rect 18170 22750 18180 22910
rect 18120 22730 18180 22750
rect 18230 22910 18290 23270
rect 18230 22750 18240 22910
rect 18280 22750 18290 22910
rect 18230 22730 18290 22750
rect 18340 22910 18400 22930
rect 18340 22750 18350 22910
rect 18390 22750 18400 22910
rect 18340 22730 18400 22750
rect 18450 22910 18510 23270
rect 18450 22750 18460 22910
rect 18500 22750 18510 22910
rect 18450 22730 18510 22750
rect 18560 22910 18620 22930
rect 18560 22750 18570 22910
rect 18610 22750 18620 22910
rect 18560 22730 18620 22750
rect 18670 22910 18730 23270
rect 18670 22750 18680 22910
rect 18720 22750 18730 22910
rect 18670 22730 18730 22750
rect 18780 22910 18840 22930
rect 18780 22750 18790 22910
rect 18830 22750 18840 22910
rect 18780 22730 18840 22750
rect 18890 22910 18950 23270
rect 18890 22750 18900 22910
rect 18940 22750 18950 22910
rect 18890 22730 18950 22750
rect 19000 22910 19060 22930
rect 19000 22750 19010 22910
rect 19050 22750 19060 22910
rect 19000 22730 19060 22750
rect 19110 22910 19170 23270
rect 19110 22750 19120 22910
rect 19160 22750 19170 22910
rect 19110 22730 19170 22750
rect 19220 22910 19280 22930
rect 19220 22750 19230 22910
rect 19270 22750 19280 22910
rect 19220 22730 19280 22750
rect 19330 22910 19390 23270
rect 19330 22750 19340 22910
rect 19380 22750 19390 22910
rect 19330 22730 19390 22750
rect 19440 22910 19500 22930
rect 19440 22750 19450 22910
rect 19490 22750 19500 22910
rect 19440 22730 19500 22750
rect 19550 22910 19610 23270
rect 19550 22750 19560 22910
rect 19600 22750 19610 22910
rect 19550 22730 19610 22750
rect 19660 22910 19720 22930
rect 19660 22750 19670 22910
rect 19710 22750 19720 22910
rect 19660 22730 19720 22750
rect 19770 22910 19830 23270
rect 19770 22750 19780 22910
rect 19820 22750 19830 22910
rect 19770 22730 19830 22750
rect 19880 22910 19940 22930
rect 19880 22750 19890 22910
rect 19930 22750 19940 22910
rect 19880 22730 19940 22750
rect 19990 22910 20050 23270
rect 19990 22750 20000 22910
rect 20040 22750 20050 22910
rect 19990 22730 20050 22750
rect 20100 22910 20160 22930
rect 20100 22750 20110 22910
rect 20150 22750 20160 22910
rect 20100 22730 20160 22750
rect 20210 22910 20270 23270
rect 20210 22750 20220 22910
rect 20260 22750 20270 22910
rect 20210 22730 20270 22750
rect 20320 22910 20380 22930
rect 20320 22750 20330 22910
rect 20370 22750 20380 22910
rect 20320 22730 20380 22750
rect 20430 22910 20490 23270
rect 20430 22750 20440 22910
rect 20480 22750 20490 22910
rect 20430 22730 20490 22750
rect 20540 22910 20600 22930
rect 20540 22750 20550 22910
rect 20590 22750 20600 22910
rect 20540 22690 20600 22750
rect 14890 22630 14900 22670
rect 14940 22630 14950 22670
rect 14110 22550 14190 22560
rect 14110 22510 14130 22550
rect 14170 22510 14190 22550
rect 14110 22500 14190 22510
rect 14330 22550 14410 22560
rect 14330 22510 14350 22550
rect 14390 22510 14410 22550
rect 14330 22500 14410 22510
rect 14550 22550 14630 22560
rect 14550 22510 14570 22550
rect 14610 22510 14630 22550
rect 14550 22500 14630 22510
rect 14770 22550 14850 22560
rect 14770 22510 14790 22550
rect 14830 22510 14850 22550
rect 14770 22500 14850 22510
rect 14110 21660 14190 21670
rect 14110 21620 14130 21660
rect 14170 21620 14190 21660
rect 14110 21610 14190 21620
rect 14330 21660 14410 21670
rect 14330 21620 14350 21660
rect 14390 21620 14410 21660
rect 14330 21610 14410 21620
rect 14550 21660 14630 21670
rect 14550 21620 14570 21660
rect 14610 21620 14630 21660
rect 14550 21610 14630 21620
rect 14770 21660 14850 21670
rect 14770 21620 14790 21660
rect 14830 21620 14850 21660
rect 14770 21610 14850 21620
rect 13890 21090 13900 21550
rect 13940 21090 13950 21550
rect 13890 21070 13950 21090
rect 14010 21550 14070 21570
rect 14010 21090 14020 21550
rect 14060 21090 14070 21550
rect 14010 21070 14070 21090
rect 14120 21550 14180 21570
rect 14120 21090 14130 21550
rect 14170 21090 14180 21550
rect 14120 21010 14180 21090
rect 14230 21550 14290 21570
rect 14230 21090 14240 21550
rect 14280 21090 14290 21550
rect 14230 21070 14290 21090
rect 14340 21550 14400 21570
rect 14340 21090 14350 21550
rect 14390 21090 14400 21550
rect 14340 21010 14400 21090
rect 14450 21550 14510 21570
rect 14450 21090 14460 21550
rect 14500 21090 14510 21550
rect 14450 21070 14510 21090
rect 14560 21550 14620 21570
rect 14560 21090 14570 21550
rect 14610 21090 14620 21550
rect 14560 21010 14620 21090
rect 14670 21550 14730 21570
rect 14670 21090 14680 21550
rect 14720 21090 14730 21550
rect 14670 21070 14730 21090
rect 14780 21550 14840 21570
rect 14780 21090 14790 21550
rect 14830 21090 14840 21550
rect 14780 21010 14840 21090
rect 14890 21550 14950 22630
rect 15080 22670 15140 22690
rect 15080 22630 15090 22670
rect 15130 22630 15140 22670
rect 15080 22610 15140 22630
rect 16830 22680 16960 22690
rect 16830 22630 16890 22680
rect 16940 22630 16960 22680
rect 16830 22620 16960 22630
rect 17020 22670 17090 22690
rect 17020 22630 17040 22670
rect 17080 22630 17090 22670
rect 15170 22550 15250 22560
rect 15170 22510 15190 22550
rect 15230 22510 15250 22550
rect 15170 22500 15250 22510
rect 15390 22550 15470 22560
rect 15390 22510 15410 22550
rect 15450 22510 15470 22550
rect 15390 22500 15470 22510
rect 15610 22550 15690 22560
rect 15610 22510 15630 22550
rect 15670 22510 15690 22550
rect 15610 22500 15690 22510
rect 15830 22550 15910 22560
rect 15830 22510 15850 22550
rect 15890 22510 15910 22550
rect 15830 22500 15910 22510
rect 16050 22550 16130 22560
rect 16050 22510 16070 22550
rect 16110 22510 16130 22550
rect 16050 22500 16130 22510
rect 16270 22550 16350 22560
rect 16270 22510 16290 22550
rect 16330 22510 16350 22550
rect 16270 22500 16350 22510
rect 16490 22550 16570 22560
rect 16490 22510 16510 22550
rect 16550 22510 16570 22550
rect 16490 22500 16570 22510
rect 16710 22550 16790 22560
rect 16710 22510 16730 22550
rect 16770 22510 16790 22550
rect 16710 22500 16790 22510
rect 15170 21660 15250 21670
rect 15170 21620 15190 21660
rect 15230 21620 15250 21660
rect 15170 21610 15250 21620
rect 15390 21660 15470 21670
rect 15390 21620 15410 21660
rect 15450 21620 15470 21660
rect 15390 21610 15470 21620
rect 15610 21660 15690 21670
rect 15610 21620 15630 21660
rect 15670 21620 15690 21660
rect 15610 21610 15690 21620
rect 15830 21660 15910 21670
rect 15830 21620 15850 21660
rect 15890 21620 15910 21660
rect 15830 21610 15910 21620
rect 16050 21660 16130 21670
rect 16050 21620 16070 21660
rect 16110 21620 16130 21660
rect 16050 21610 16130 21620
rect 16270 21660 16350 21670
rect 16270 21620 16290 21660
rect 16330 21620 16350 21660
rect 16270 21610 16350 21620
rect 16490 21660 16570 21670
rect 16490 21620 16510 21660
rect 16550 21620 16570 21660
rect 16490 21610 16570 21620
rect 16710 21660 16790 21670
rect 16710 21620 16730 21660
rect 16770 21620 16790 21660
rect 16710 21610 16790 21620
rect 14890 21090 14900 21550
rect 14940 21090 14950 21550
rect 14890 21070 14950 21090
rect 15070 21550 15130 21570
rect 15070 21090 15080 21550
rect 15120 21090 15130 21550
rect 15070 21070 15130 21090
rect 15180 21550 15240 21570
rect 15180 21090 15190 21550
rect 15230 21090 15240 21550
rect 15180 21010 15240 21090
rect 15290 21550 15350 21570
rect 15290 21090 15300 21550
rect 15340 21090 15350 21550
rect 15290 21070 15350 21090
rect 15400 21550 15460 21570
rect 15400 21090 15410 21550
rect 15450 21090 15460 21550
rect 15400 21010 15460 21090
rect 15510 21550 15570 21570
rect 15510 21090 15520 21550
rect 15560 21090 15570 21550
rect 15510 21070 15570 21090
rect 15620 21550 15680 21570
rect 15620 21090 15630 21550
rect 15670 21090 15680 21550
rect 15620 21010 15680 21090
rect 15730 21550 15790 21570
rect 15730 21090 15740 21550
rect 15780 21090 15790 21550
rect 15730 21070 15790 21090
rect 15840 21550 15900 21570
rect 15840 21090 15850 21550
rect 15890 21090 15900 21550
rect 15840 21010 15900 21090
rect 15950 21550 16010 21570
rect 15950 21090 15960 21550
rect 16000 21090 16010 21550
rect 15950 21070 16010 21090
rect 16060 21550 16120 21570
rect 16060 21090 16070 21550
rect 16110 21090 16120 21550
rect 16060 21010 16120 21090
rect 16170 21550 16230 21570
rect 16170 21090 16180 21550
rect 16220 21090 16230 21550
rect 16170 21070 16230 21090
rect 16280 21550 16340 21570
rect 16280 21090 16290 21550
rect 16330 21090 16340 21550
rect 16280 21010 16340 21090
rect 16390 21550 16450 21570
rect 16390 21090 16400 21550
rect 16440 21090 16450 21550
rect 16390 21070 16450 21090
rect 16500 21550 16560 21570
rect 16500 21090 16510 21550
rect 16550 21090 16560 21550
rect 16500 21010 16560 21090
rect 16610 21550 16670 21570
rect 16610 21090 16620 21550
rect 16660 21090 16670 21550
rect 16610 21070 16670 21090
rect 16720 21550 16780 21570
rect 16720 21090 16730 21550
rect 16770 21090 16780 21550
rect 16720 21010 16780 21090
rect 16830 21550 16890 22620
rect 17020 22610 17090 22630
rect 20540 22680 20670 22690
rect 20540 22630 20600 22680
rect 20650 22630 20670 22680
rect 20540 22620 20670 22630
rect 17120 22550 17200 22560
rect 17120 22510 17140 22550
rect 17180 22510 17200 22550
rect 17120 22500 17200 22510
rect 17340 22550 17420 22560
rect 17340 22510 17360 22550
rect 17400 22510 17420 22550
rect 17340 22500 17420 22510
rect 17560 22550 17640 22560
rect 17560 22510 17580 22550
rect 17620 22510 17640 22550
rect 17560 22500 17640 22510
rect 17780 22550 17860 22560
rect 17780 22510 17800 22550
rect 17840 22510 17860 22550
rect 17780 22500 17860 22510
rect 18000 22550 18080 22560
rect 18000 22510 18020 22550
rect 18060 22510 18080 22550
rect 18000 22500 18080 22510
rect 18220 22550 18300 22560
rect 18220 22510 18240 22550
rect 18280 22510 18300 22550
rect 18220 22500 18300 22510
rect 18440 22550 18520 22560
rect 18440 22510 18460 22550
rect 18500 22510 18520 22550
rect 18440 22500 18520 22510
rect 18660 22550 18740 22560
rect 18660 22510 18680 22550
rect 18720 22510 18740 22550
rect 18660 22500 18740 22510
rect 18880 22550 18960 22560
rect 18880 22510 18900 22550
rect 18940 22510 18960 22550
rect 18880 22500 18960 22510
rect 19100 22550 19180 22560
rect 19100 22510 19120 22550
rect 19160 22510 19180 22550
rect 19100 22500 19180 22510
rect 19320 22550 19400 22560
rect 19320 22510 19340 22550
rect 19380 22510 19400 22550
rect 19320 22500 19400 22510
rect 19540 22550 19620 22560
rect 19540 22510 19560 22550
rect 19600 22510 19620 22550
rect 19540 22500 19620 22510
rect 19760 22550 19840 22560
rect 19760 22510 19780 22550
rect 19820 22510 19840 22550
rect 19760 22500 19840 22510
rect 19980 22550 20060 22560
rect 19980 22510 20000 22550
rect 20040 22510 20060 22550
rect 19980 22500 20060 22510
rect 20200 22550 20280 22560
rect 20200 22510 20220 22550
rect 20260 22510 20280 22550
rect 20200 22500 20280 22510
rect 20420 22550 20500 22560
rect 20420 22510 20440 22550
rect 20480 22510 20500 22550
rect 20420 22500 20500 22510
rect 17120 21660 17200 21670
rect 17120 21620 17140 21660
rect 17180 21620 17200 21660
rect 17120 21610 17200 21620
rect 17340 21660 17420 21670
rect 17340 21620 17360 21660
rect 17400 21620 17420 21660
rect 17340 21610 17420 21620
rect 17560 21660 17640 21670
rect 17560 21620 17580 21660
rect 17620 21620 17640 21660
rect 17560 21610 17640 21620
rect 17780 21660 17860 21670
rect 17780 21620 17800 21660
rect 17840 21620 17860 21660
rect 17780 21610 17860 21620
rect 18000 21660 18080 21670
rect 18000 21620 18020 21660
rect 18060 21620 18080 21660
rect 18000 21610 18080 21620
rect 18220 21660 18300 21670
rect 18220 21620 18240 21660
rect 18280 21620 18300 21660
rect 18220 21610 18300 21620
rect 18440 21660 18520 21670
rect 18440 21620 18460 21660
rect 18500 21620 18520 21660
rect 18440 21610 18520 21620
rect 18660 21660 18740 21670
rect 18660 21620 18680 21660
rect 18720 21620 18740 21660
rect 18660 21610 18740 21620
rect 18880 21660 18960 21670
rect 18880 21620 18900 21660
rect 18940 21620 18960 21660
rect 18880 21610 18960 21620
rect 19100 21660 19180 21670
rect 19100 21620 19120 21660
rect 19160 21620 19180 21660
rect 19100 21610 19180 21620
rect 19320 21660 19400 21670
rect 19320 21620 19340 21660
rect 19380 21620 19400 21660
rect 19320 21610 19400 21620
rect 19540 21660 19620 21670
rect 19540 21620 19560 21660
rect 19600 21620 19620 21660
rect 19540 21610 19620 21620
rect 19760 21660 19840 21670
rect 19760 21620 19780 21660
rect 19820 21620 19840 21660
rect 19760 21610 19840 21620
rect 19980 21660 20060 21670
rect 19980 21620 20000 21660
rect 20040 21620 20060 21660
rect 19980 21610 20060 21620
rect 20200 21660 20280 21670
rect 20200 21620 20220 21660
rect 20260 21620 20280 21660
rect 20200 21610 20280 21620
rect 20420 21660 20500 21670
rect 20420 21620 20440 21660
rect 20480 21620 20500 21660
rect 20420 21610 20500 21620
rect 16830 21090 16840 21550
rect 16880 21090 16890 21550
rect 16830 21070 16890 21090
rect 17020 21550 17080 21570
rect 17020 21090 17030 21550
rect 17070 21090 17080 21550
rect 17020 21070 17080 21090
rect 17130 21550 17190 21570
rect 17130 21090 17140 21550
rect 17180 21090 17190 21550
rect 17130 21010 17190 21090
rect 17240 21550 17300 21570
rect 17240 21090 17250 21550
rect 17290 21090 17300 21550
rect 17240 21070 17300 21090
rect 17350 21550 17410 21570
rect 17350 21090 17360 21550
rect 17400 21090 17410 21550
rect 17350 21010 17410 21090
rect 17460 21550 17520 21570
rect 17460 21090 17470 21550
rect 17510 21090 17520 21550
rect 17460 21070 17520 21090
rect 17570 21550 17630 21570
rect 17570 21090 17580 21550
rect 17620 21090 17630 21550
rect 17570 21010 17630 21090
rect 17680 21550 17740 21570
rect 17680 21090 17690 21550
rect 17730 21090 17740 21550
rect 17680 21070 17740 21090
rect 17790 21550 17850 21570
rect 17790 21090 17800 21550
rect 17840 21090 17850 21550
rect 17790 21010 17850 21090
rect 17900 21550 17960 21570
rect 17900 21090 17910 21550
rect 17950 21090 17960 21550
rect 17900 21070 17960 21090
rect 18010 21550 18070 21570
rect 18010 21090 18020 21550
rect 18060 21090 18070 21550
rect 18010 21010 18070 21090
rect 18120 21550 18180 21570
rect 18120 21090 18130 21550
rect 18170 21090 18180 21550
rect 18120 21070 18180 21090
rect 18230 21550 18290 21570
rect 18230 21090 18240 21550
rect 18280 21090 18290 21550
rect 18230 21010 18290 21090
rect 18340 21550 18400 21570
rect 18340 21090 18350 21550
rect 18390 21090 18400 21550
rect 18340 21070 18400 21090
rect 18450 21550 18510 21570
rect 18450 21090 18460 21550
rect 18500 21090 18510 21550
rect 18450 21010 18510 21090
rect 18560 21550 18620 21570
rect 18560 21090 18570 21550
rect 18610 21090 18620 21550
rect 18560 21070 18620 21090
rect 18670 21550 18730 21570
rect 18670 21090 18680 21550
rect 18720 21090 18730 21550
rect 18670 21010 18730 21090
rect 18780 21550 18840 21570
rect 18780 21090 18790 21550
rect 18830 21090 18840 21550
rect 18780 21070 18840 21090
rect 18890 21550 18950 21570
rect 18890 21090 18900 21550
rect 18940 21090 18950 21550
rect 18890 21010 18950 21090
rect 19000 21550 19060 21570
rect 19000 21090 19010 21550
rect 19050 21090 19060 21550
rect 19000 21070 19060 21090
rect 19110 21550 19170 21570
rect 19110 21090 19120 21550
rect 19160 21090 19170 21550
rect 19110 21010 19170 21090
rect 19220 21550 19280 21570
rect 19220 21090 19230 21550
rect 19270 21090 19280 21550
rect 19220 21070 19280 21090
rect 19330 21550 19390 21570
rect 19330 21090 19340 21550
rect 19380 21090 19390 21550
rect 19330 21010 19390 21090
rect 19440 21550 19500 21570
rect 19440 21090 19450 21550
rect 19490 21090 19500 21550
rect 19440 21070 19500 21090
rect 19550 21550 19610 21570
rect 19550 21090 19560 21550
rect 19600 21090 19610 21550
rect 19550 21010 19610 21090
rect 19660 21550 19720 21570
rect 19660 21090 19670 21550
rect 19710 21090 19720 21550
rect 19660 21070 19720 21090
rect 19770 21550 19830 21570
rect 19770 21090 19780 21550
rect 19820 21090 19830 21550
rect 19770 21010 19830 21090
rect 19880 21550 19940 21570
rect 19880 21090 19890 21550
rect 19930 21090 19940 21550
rect 19880 21070 19940 21090
rect 19990 21550 20050 21570
rect 19990 21090 20000 21550
rect 20040 21090 20050 21550
rect 19990 21010 20050 21090
rect 20100 21550 20160 21570
rect 20100 21090 20110 21550
rect 20150 21090 20160 21550
rect 20100 21070 20160 21090
rect 20210 21550 20270 21570
rect 20210 21090 20220 21550
rect 20260 21090 20270 21550
rect 20210 21010 20270 21090
rect 20320 21550 20380 21570
rect 20320 21090 20330 21550
rect 20370 21090 20380 21550
rect 20320 21070 20380 21090
rect 20430 21550 20490 21570
rect 20430 21090 20440 21550
rect 20480 21090 20490 21550
rect 20430 21010 20490 21090
rect 20540 21550 20600 22620
rect 20540 21090 20550 21550
rect 20590 21090 20600 21550
rect 20540 21070 20600 21090
rect 7280 21000 20640 21010
rect 7280 20960 7320 21000
rect 7360 20960 7400 21000
rect 7440 20960 7480 21000
rect 7520 20960 7560 21000
rect 7600 20960 7640 21000
rect 7680 20960 7720 21000
rect 7760 20960 7800 21000
rect 7840 20960 7880 21000
rect 7920 20960 7960 21000
rect 8000 20960 8040 21000
rect 8080 20960 8120 21000
rect 8160 20960 8200 21000
rect 8240 20960 8280 21000
rect 8320 20960 8360 21000
rect 8400 20960 8440 21000
rect 8480 20960 8520 21000
rect 8560 20960 8600 21000
rect 8640 20960 8680 21000
rect 8720 20960 8760 21000
rect 8800 20960 8840 21000
rect 8880 20960 8920 21000
rect 8960 20960 9000 21000
rect 9040 20960 9080 21000
rect 9120 20960 9160 21000
rect 9200 20960 9260 21000
rect 9300 20960 9340 21000
rect 9380 20960 9420 21000
rect 9460 20960 9500 21000
rect 9540 20960 9580 21000
rect 9620 20960 9660 21000
rect 9700 20960 9740 21000
rect 9780 20960 9820 21000
rect 9860 20960 9900 21000
rect 9940 20960 9980 21000
rect 10020 20960 10060 21000
rect 10100 20960 10140 21000
rect 10180 20960 10220 21000
rect 10260 20960 10300 21000
rect 10340 20960 10380 21000
rect 10420 20960 10460 21000
rect 10500 20960 10540 21000
rect 10580 20960 10620 21000
rect 10660 20960 10700 21000
rect 10740 20960 10780 21000
rect 10820 20960 10860 21000
rect 10900 20960 10940 21000
rect 10980 20960 11020 21000
rect 11060 20960 11100 21000
rect 11140 20960 11180 21000
rect 11220 20960 11260 21000
rect 11300 20960 11340 21000
rect 11380 20960 11420 21000
rect 11460 20960 11500 21000
rect 11540 20960 11580 21000
rect 11620 20960 11660 21000
rect 11700 20960 11740 21000
rect 11780 20960 11820 21000
rect 11860 20960 11900 21000
rect 11940 20960 11980 21000
rect 12020 20960 12060 21000
rect 12100 20960 12140 21000
rect 12180 20960 12220 21000
rect 12260 20960 12300 21000
rect 12340 20960 12380 21000
rect 12420 20960 12460 21000
rect 12500 20960 12540 21000
rect 12580 20960 12620 21000
rect 12660 20960 12700 21000
rect 12740 20960 12780 21000
rect 12820 20960 12880 21000
rect 12920 20960 12960 21000
rect 13000 20960 13040 21000
rect 13080 20960 13120 21000
rect 13160 20960 13200 21000
rect 13240 20960 13280 21000
rect 13320 20960 13360 21000
rect 13400 20960 13440 21000
rect 13480 20960 13520 21000
rect 13560 20960 13600 21000
rect 13640 20960 13680 21000
rect 13720 20960 13760 21000
rect 13800 20960 13840 21000
rect 13880 20960 13920 21000
rect 13960 20960 14000 21000
rect 14040 20960 14080 21000
rect 14120 20960 14160 21000
rect 14200 20960 14240 21000
rect 14280 20960 14320 21000
rect 14360 20960 14400 21000
rect 14440 20960 14480 21000
rect 14520 20960 14560 21000
rect 14600 20960 14640 21000
rect 14680 20960 14720 21000
rect 14760 20960 14800 21000
rect 14840 20960 14880 21000
rect 14920 20960 14960 21000
rect 15000 20960 15040 21000
rect 15080 20960 15120 21000
rect 15160 20960 15200 21000
rect 15240 20960 15280 21000
rect 15320 20960 15360 21000
rect 15400 20960 15440 21000
rect 15480 20960 15520 21000
rect 15560 20960 15600 21000
rect 15640 20960 15680 21000
rect 15720 20960 15760 21000
rect 15800 20960 15840 21000
rect 15880 20960 15920 21000
rect 15960 20960 16000 21000
rect 16040 20960 16080 21000
rect 16120 20960 16160 21000
rect 16200 20960 16240 21000
rect 16280 20960 16320 21000
rect 16360 20960 16400 21000
rect 16440 20960 16480 21000
rect 16520 20960 16560 21000
rect 16600 20960 16640 21000
rect 16680 20960 16720 21000
rect 16760 20960 16800 21000
rect 16840 20960 16880 21000
rect 16920 20960 16960 21000
rect 17000 20960 17040 21000
rect 17080 20960 17120 21000
rect 17160 20960 17200 21000
rect 17240 20960 17280 21000
rect 17320 20960 17360 21000
rect 17400 20960 17440 21000
rect 17480 20960 17520 21000
rect 17560 20960 17600 21000
rect 17640 20960 17680 21000
rect 17720 20960 17760 21000
rect 17800 20960 17840 21000
rect 17880 20960 17920 21000
rect 17960 20960 18000 21000
rect 18040 20960 18080 21000
rect 18120 20960 18160 21000
rect 18200 20960 18240 21000
rect 18280 20960 18320 21000
rect 18360 20960 18400 21000
rect 18440 20960 18480 21000
rect 18520 20960 18560 21000
rect 18600 20960 18640 21000
rect 18680 20960 18720 21000
rect 18760 20960 18800 21000
rect 18840 20960 18880 21000
rect 18920 20960 18960 21000
rect 19000 20960 19040 21000
rect 19080 20960 19120 21000
rect 19160 20960 19200 21000
rect 19240 20960 19280 21000
rect 19320 20960 19360 21000
rect 19400 20960 19440 21000
rect 19480 20960 19520 21000
rect 19560 20960 19600 21000
rect 19640 20960 19680 21000
rect 19720 20960 19760 21000
rect 19800 20960 19840 21000
rect 19880 20960 19920 21000
rect 19960 20960 20000 21000
rect 20040 20960 20080 21000
rect 20120 20960 20160 21000
rect 20200 20960 20240 21000
rect 20280 20960 20320 21000
rect 20360 20960 20400 21000
rect 20440 20960 20480 21000
rect 20520 20960 20560 21000
rect 20600 20960 20640 21000
rect 7280 20950 20640 20960
rect 7280 20470 8230 20480
rect 7280 20430 7320 20470
rect 7360 20430 7400 20470
rect 7440 20430 7480 20470
rect 7520 20430 7560 20470
rect 7600 20430 7640 20470
rect 7680 20430 7720 20470
rect 7760 20430 7800 20470
rect 7840 20430 7880 20470
rect 7920 20430 7960 20470
rect 8000 20430 8040 20470
rect 8080 20430 8120 20470
rect 8160 20430 8230 20470
rect 7280 20420 8230 20430
rect 7390 20340 7450 20420
rect 7390 19380 7400 20340
rect 7440 19380 7450 20340
rect 7390 19360 7450 19380
rect 7650 20340 7710 20360
rect 7650 19380 7660 20340
rect 7700 19380 7710 20340
rect 7950 20340 8010 20420
rect 7950 19880 7960 20340
rect 8000 19880 8010 20340
rect 7950 19860 8010 19880
rect 8060 20340 8120 20360
rect 8060 19880 8070 20340
rect 8110 19880 8120 20340
rect 7350 19310 7490 19320
rect 7350 19270 7400 19310
rect 7440 19270 7490 19310
rect 7350 19260 7490 19270
rect 7350 18430 7490 18440
rect 7350 18390 7400 18430
rect 7440 18390 7490 18430
rect 7350 18380 7490 18390
rect 7650 18360 7710 19380
rect 8060 18360 8120 19880
rect 8170 20340 8230 20420
rect 8170 19880 8180 20340
rect 8220 19880 8230 20340
rect 8310 20020 20640 20030
rect 8310 19980 8360 20020
rect 8400 19980 8440 20020
rect 8480 19980 8520 20020
rect 8560 19980 8600 20020
rect 8640 19980 8680 20020
rect 8720 19980 8760 20020
rect 8800 19980 8840 20020
rect 8880 19980 8920 20020
rect 8960 19980 9000 20020
rect 9040 19980 9080 20020
rect 9120 19980 9160 20020
rect 9200 19980 9260 20020
rect 9300 19980 9340 20020
rect 9380 19980 9420 20020
rect 9460 19980 9500 20020
rect 9540 19980 9580 20020
rect 9620 19980 9660 20020
rect 9700 19980 9740 20020
rect 9780 19980 9820 20020
rect 9860 19980 9900 20020
rect 9940 19980 9980 20020
rect 10020 19980 10060 20020
rect 10100 19980 10140 20020
rect 10180 19980 10220 20020
rect 10260 19980 10300 20020
rect 10340 19980 10380 20020
rect 10420 19980 10460 20020
rect 10500 19980 10540 20020
rect 10580 19980 10620 20020
rect 10660 19980 10700 20020
rect 10740 19980 10780 20020
rect 10820 19980 10860 20020
rect 10900 19980 10940 20020
rect 10980 19980 11020 20020
rect 11060 19980 11100 20020
rect 11140 19980 11180 20020
rect 11220 19980 11260 20020
rect 11300 19980 11340 20020
rect 11380 19980 11420 20020
rect 11460 19980 11500 20020
rect 11540 19980 11580 20020
rect 11620 19980 11660 20020
rect 11700 19980 11740 20020
rect 11780 19980 11820 20020
rect 11860 19980 11900 20020
rect 11940 19980 11980 20020
rect 12020 19980 12060 20020
rect 12100 19980 12140 20020
rect 12180 19980 12220 20020
rect 12260 19980 12300 20020
rect 12340 19980 12380 20020
rect 12420 19980 12460 20020
rect 12500 19980 12540 20020
rect 12580 19980 12620 20020
rect 12660 19980 12700 20020
rect 12740 19980 12780 20020
rect 12820 19980 12860 20020
rect 12900 19980 12940 20020
rect 12980 19980 13040 20020
rect 13080 19980 13120 20020
rect 13160 19980 13200 20020
rect 13240 19980 13280 20020
rect 13320 19980 13360 20020
rect 13400 19980 13440 20020
rect 13480 19980 13520 20020
rect 13560 19980 13600 20020
rect 13640 19980 13680 20020
rect 13720 19980 13760 20020
rect 13800 19980 13840 20020
rect 13880 19980 13920 20020
rect 13960 19980 14000 20020
rect 14040 19980 14080 20020
rect 14120 19980 14160 20020
rect 14200 19980 14240 20020
rect 14280 19980 14320 20020
rect 14360 19980 14400 20020
rect 14440 19980 14480 20020
rect 14520 19980 14560 20020
rect 14600 19980 14640 20020
rect 14680 19980 14720 20020
rect 14760 19980 14800 20020
rect 14840 19980 14880 20020
rect 14920 19980 14960 20020
rect 15000 19980 15040 20020
rect 15080 19980 15120 20020
rect 15160 19980 15200 20020
rect 15240 19980 15280 20020
rect 15320 19980 15360 20020
rect 15400 19980 15440 20020
rect 15480 19980 15520 20020
rect 15560 19980 15600 20020
rect 15640 19980 15680 20020
rect 15720 19980 15760 20020
rect 15800 19980 15840 20020
rect 15880 19980 15920 20020
rect 15960 19980 16000 20020
rect 16040 19980 16080 20020
rect 16120 19980 16160 20020
rect 16200 19980 16240 20020
rect 16280 19980 16320 20020
rect 16360 19980 16400 20020
rect 16440 19980 16480 20020
rect 16520 19980 16560 20020
rect 16600 19980 16640 20020
rect 16680 19980 16720 20020
rect 16760 19980 16800 20020
rect 16840 19980 16880 20020
rect 16920 19980 16960 20020
rect 17000 19980 17040 20020
rect 17080 19980 17120 20020
rect 17160 19980 17200 20020
rect 17240 19980 17280 20020
rect 17320 19980 17360 20020
rect 17400 19980 17440 20020
rect 17480 19980 17520 20020
rect 17560 19980 17600 20020
rect 17640 19980 17680 20020
rect 17720 19980 17760 20020
rect 17800 19980 17840 20020
rect 17880 19980 17920 20020
rect 17960 19980 18000 20020
rect 18040 19980 18080 20020
rect 18120 19980 18160 20020
rect 18200 19980 18240 20020
rect 18280 19980 18320 20020
rect 18360 19980 18400 20020
rect 18440 19980 18480 20020
rect 18520 19980 18560 20020
rect 18600 19980 18640 20020
rect 18680 19980 18720 20020
rect 18760 19980 18800 20020
rect 18840 19980 18880 20020
rect 18920 19980 18960 20020
rect 19000 19980 19040 20020
rect 19080 19980 19120 20020
rect 19160 19980 19200 20020
rect 19240 19980 19280 20020
rect 19320 19980 19360 20020
rect 19400 19980 19440 20020
rect 19480 19980 19520 20020
rect 19560 19980 19600 20020
rect 19640 19980 19680 20020
rect 19720 19980 19760 20020
rect 19800 19980 19840 20020
rect 19880 19980 19920 20020
rect 19960 19980 20000 20020
rect 20040 19980 20080 20020
rect 20120 19980 20160 20020
rect 20200 19980 20240 20020
rect 20280 19980 20320 20020
rect 20360 19980 20400 20020
rect 20440 19980 20480 20020
rect 20520 19980 20560 20020
rect 20600 19980 20640 20020
rect 8310 19970 20640 19980
rect 8170 19860 8230 19880
rect 8480 19890 8540 19970
rect 8480 19430 8490 19890
rect 8530 19430 8540 19890
rect 8480 19410 8540 19430
rect 8610 19890 8670 19910
rect 8610 19430 8620 19890
rect 8660 19430 8670 19890
rect 8610 18370 8670 19430
rect 8740 19890 8800 19970
rect 8740 19430 8750 19890
rect 8790 19430 8800 19890
rect 8740 19410 8800 19430
rect 8860 19890 8920 19970
rect 8860 19430 8870 19890
rect 8910 19430 8920 19890
rect 8860 19410 8920 19430
rect 8970 19890 9030 19910
rect 8970 19430 8980 19890
rect 9020 19430 9030 19890
rect 8970 18370 9030 19430
rect 9220 19890 9280 19970
rect 9220 19430 9230 19890
rect 9270 19430 9280 19890
rect 9220 19410 9280 19430
rect 9330 19890 9390 19910
rect 9330 19430 9340 19890
rect 9380 19430 9390 19890
rect 7650 18300 7820 18360
rect 8060 18300 8230 18360
rect 7550 18280 7610 18300
rect 7550 18240 7560 18280
rect 7600 18240 7610 18280
rect 7550 18220 7610 18240
rect 7290 18170 7350 18190
rect 7290 18130 7300 18170
rect 7340 18130 7350 18170
rect 7290 18110 7350 18130
rect 7760 18070 7820 18300
rect 7960 18280 8020 18300
rect 7960 18240 7970 18280
rect 8010 18240 8020 18280
rect 7960 18220 8020 18240
rect 8170 18080 8230 18300
rect 8480 18350 8550 18370
rect 8480 18310 8500 18350
rect 8540 18310 8550 18350
rect 8610 18350 8930 18370
rect 8610 18330 8800 18350
rect 8480 18290 8550 18310
rect 8740 18310 8800 18330
rect 8840 18310 8880 18350
rect 8920 18310 8930 18350
rect 8740 18290 8930 18310
rect 8970 18350 9160 18370
rect 8970 18310 9000 18350
rect 9040 18310 9160 18350
rect 8970 18290 9160 18310
rect 8630 18270 8700 18290
rect 8630 18230 8650 18270
rect 8690 18230 8700 18270
rect 8630 18210 8700 18230
rect 7280 18030 7780 18070
rect 7280 18020 7820 18030
rect 7280 17960 7340 18020
rect 7280 17800 7290 17960
rect 7330 17800 7340 17960
rect 7280 17780 7340 17800
rect 7390 17960 7450 17980
rect 7390 17800 7400 17960
rect 7440 17800 7450 17960
rect 7390 17710 7450 17800
rect 7520 17960 7580 18020
rect 7520 17800 7530 17960
rect 7570 17800 7580 17960
rect 7520 17780 7580 17800
rect 7650 17960 7710 17980
rect 7650 17800 7660 17960
rect 7700 17800 7710 17960
rect 7650 17710 7710 17800
rect 7760 17960 7820 18020
rect 8060 18070 8230 18080
rect 8060 18030 8190 18070
rect 8060 18020 8230 18030
rect 8480 18150 8540 18170
rect 7760 17800 7770 17960
rect 7810 17800 7820 17960
rect 7760 17780 7820 17800
rect 7950 17960 8010 17980
rect 7950 17800 7960 17960
rect 8000 17800 8010 17960
rect 7950 17710 8010 17800
rect 8060 17960 8120 18020
rect 8060 17800 8070 17960
rect 8110 17800 8120 17960
rect 8060 17780 8120 17800
rect 8170 17960 8230 17980
rect 8170 17800 8180 17960
rect 8220 17800 8230 17960
rect 8170 17710 8230 17800
rect 8480 17790 8490 18150
rect 8530 17790 8540 18150
rect 8480 17710 8540 17790
rect 8610 18150 8670 18170
rect 8610 17790 8620 18150
rect 8660 17790 8670 18150
rect 8610 17770 8670 17790
rect 8740 18150 8800 18290
rect 8740 17790 8750 18150
rect 8790 17790 8800 18150
rect 8740 17770 8800 17790
rect 8860 18220 8920 18240
rect 8860 18060 8870 18220
rect 8910 18060 8920 18220
rect 8860 17710 8920 18060
rect 8970 18220 9030 18290
rect 8970 18060 8980 18220
rect 9020 18060 9030 18220
rect 9090 18200 9160 18290
rect 9200 18330 9290 18350
rect 9200 18270 9220 18330
rect 9280 18270 9290 18330
rect 9200 18250 9290 18270
rect 9330 18250 9390 19430
rect 9440 19890 9500 19970
rect 9440 19430 9450 19890
rect 9490 19430 9500 19890
rect 9440 19410 9500 19430
rect 9670 19890 9730 19970
rect 9670 19430 9680 19890
rect 9720 19430 9730 19890
rect 9670 19410 9730 19430
rect 9800 19890 9860 19910
rect 9800 19430 9810 19890
rect 9850 19430 9860 19890
rect 9660 19360 9740 19370
rect 9660 19320 9680 19360
rect 9720 19320 9740 19360
rect 9660 19310 9740 19320
rect 9660 18470 9740 18480
rect 9660 18430 9680 18470
rect 9720 18430 9740 18470
rect 9660 18420 9740 18430
rect 9800 18370 9860 19430
rect 9930 19890 9990 19970
rect 9930 19430 9940 19890
rect 9980 19430 9990 19890
rect 9930 19410 9990 19430
rect 10160 19890 10220 19970
rect 10160 19430 10170 19890
rect 10210 19430 10220 19890
rect 10160 19410 10220 19430
rect 10270 19890 10330 19910
rect 10270 19430 10280 19890
rect 10320 19430 10330 19890
rect 9920 19360 10000 19370
rect 9920 19320 9940 19360
rect 9980 19320 10000 19360
rect 9920 19310 10000 19320
rect 9920 18470 10000 18480
rect 9920 18430 9940 18470
rect 9980 18430 10000 18470
rect 9920 18420 10000 18430
rect 10270 18370 10330 19430
rect 10380 19890 10440 19970
rect 10380 19430 10390 19890
rect 10430 19430 10440 19890
rect 10380 19410 10440 19430
rect 10660 19890 10720 19970
rect 10660 19430 10670 19890
rect 10710 19430 10720 19890
rect 10660 19410 10720 19430
rect 10790 19890 10850 19910
rect 10790 19430 10800 19890
rect 10840 19430 10850 19890
rect 10650 19360 10730 19370
rect 10650 19320 10670 19360
rect 10710 19320 10730 19360
rect 10650 19310 10730 19320
rect 10650 18470 10730 18480
rect 10650 18430 10670 18470
rect 10710 18430 10730 18470
rect 10650 18420 10730 18430
rect 10790 18370 10850 19430
rect 10920 19890 10980 19970
rect 10920 19430 10930 19890
rect 10970 19430 10980 19890
rect 10920 19410 10980 19430
rect 11150 19890 11210 19970
rect 11150 19430 11160 19890
rect 11200 19430 11210 19890
rect 11150 19410 11210 19430
rect 11260 19890 11320 19910
rect 11260 19430 11270 19890
rect 11310 19430 11320 19890
rect 10910 19360 10990 19370
rect 10910 19320 10930 19360
rect 10970 19320 10990 19360
rect 10910 19310 10990 19320
rect 10910 18470 10990 18480
rect 10910 18430 10930 18470
rect 10970 18430 10990 18470
rect 10910 18420 10990 18430
rect 11260 18370 11320 19430
rect 11370 19890 11430 19970
rect 11370 19430 11380 19890
rect 11420 19430 11430 19890
rect 11370 19410 11430 19430
rect 11660 19890 11720 19970
rect 11660 19430 11670 19890
rect 11710 19430 11720 19890
rect 11660 19410 11720 19430
rect 11790 19890 11850 19910
rect 11790 19430 11800 19890
rect 11840 19430 11850 19890
rect 11650 19350 11730 19360
rect 11650 19310 11670 19350
rect 11710 19310 11730 19350
rect 11650 19300 11730 19310
rect 11650 18460 11730 18470
rect 11650 18420 11670 18460
rect 11710 18420 11730 18460
rect 11650 18410 11730 18420
rect 11790 18370 11850 19430
rect 11920 19890 11980 19970
rect 11920 19430 11930 19890
rect 11970 19430 11980 19890
rect 11920 19410 11980 19430
rect 12150 19890 12210 19970
rect 12150 19430 12160 19890
rect 12200 19430 12210 19890
rect 12150 19410 12210 19430
rect 12260 19890 12320 19910
rect 12260 19430 12270 19890
rect 12310 19430 12320 19890
rect 11910 19350 11990 19360
rect 11910 19310 11930 19350
rect 11970 19310 11990 19350
rect 11910 19300 11990 19310
rect 11910 18460 11990 18470
rect 11910 18420 11930 18460
rect 11970 18420 11990 18460
rect 11910 18410 11990 18420
rect 12260 18370 12320 19430
rect 12370 19890 12430 19970
rect 12370 19430 12380 19890
rect 12420 19430 12430 19890
rect 12370 19410 12430 19430
rect 12530 19890 12590 19970
rect 12530 19430 12540 19890
rect 12580 19430 12590 19890
rect 12530 19410 12590 19430
rect 12640 19890 12700 19910
rect 12640 19430 12650 19890
rect 12690 19430 12700 19890
rect 12640 18370 12700 19430
rect 12750 19890 12810 19970
rect 12750 19430 12760 19890
rect 12800 19430 12810 19890
rect 12750 19410 12810 19430
rect 12880 19890 12940 19970
rect 12880 19430 12890 19890
rect 12930 19430 12940 19890
rect 12880 19410 12940 19430
rect 12990 19890 13050 19910
rect 12990 19430 13000 19890
rect 13040 19430 13050 19890
rect 9570 18350 9630 18370
rect 9570 18310 9580 18350
rect 9620 18310 9630 18350
rect 9800 18360 10230 18370
rect 9800 18320 10080 18360
rect 10120 18320 10160 18360
rect 10200 18320 10230 18360
rect 9800 18310 10230 18320
rect 10270 18360 10510 18370
rect 10270 18320 10460 18360
rect 10500 18320 10510 18360
rect 10270 18310 10510 18320
rect 10560 18350 10620 18370
rect 10560 18310 10570 18350
rect 10610 18310 10620 18350
rect 10790 18360 11220 18370
rect 10790 18320 11070 18360
rect 11110 18320 11150 18360
rect 11190 18320 11220 18360
rect 10790 18310 11220 18320
rect 11260 18360 11500 18370
rect 11260 18320 11450 18360
rect 11490 18320 11500 18360
rect 11260 18310 11500 18320
rect 11560 18350 11620 18370
rect 11560 18310 11570 18350
rect 11610 18310 11620 18350
rect 11790 18360 12220 18370
rect 11790 18320 12070 18360
rect 12110 18320 12150 18360
rect 12190 18320 12220 18360
rect 11790 18310 12220 18320
rect 12260 18360 12600 18370
rect 12260 18320 12450 18360
rect 12490 18320 12530 18360
rect 12570 18320 12600 18360
rect 12260 18310 12600 18320
rect 12640 18350 12950 18370
rect 12640 18310 12820 18350
rect 12860 18310 12900 18350
rect 12940 18310 12950 18350
rect 9570 18290 9630 18310
rect 9830 18250 9890 18270
rect 9330 18210 9840 18250
rect 9880 18210 9890 18250
rect 9080 18180 9170 18200
rect 9080 18130 9100 18180
rect 9150 18130 9170 18180
rect 9080 18110 9170 18130
rect 8970 18040 9030 18060
rect 9220 17950 9280 17970
rect 9220 17790 9230 17950
rect 9270 17790 9280 17950
rect 9220 17710 9280 17790
rect 9330 17950 9390 18210
rect 9830 18190 9890 18210
rect 9670 18150 9730 18170
rect 9330 17790 9340 17950
rect 9380 17790 9390 17950
rect 9330 17770 9390 17790
rect 9440 17950 9500 17970
rect 9440 17790 9450 17950
rect 9490 17790 9500 17950
rect 9440 17710 9500 17790
rect 9670 17790 9680 18150
rect 9720 17790 9730 18150
rect 9670 17710 9730 17790
rect 9930 18150 9990 18310
rect 9930 17790 9940 18150
rect 9980 17790 9990 18150
rect 9930 17770 9990 17790
rect 10160 17950 10220 17970
rect 10160 17790 10170 17950
rect 10210 17790 10220 17950
rect 10160 17710 10220 17790
rect 10270 17950 10330 18310
rect 10560 18290 10620 18310
rect 10820 18250 10880 18270
rect 10820 18210 10830 18250
rect 10870 18210 10880 18250
rect 10820 18190 10880 18210
rect 10660 18150 10720 18170
rect 10270 17790 10280 17950
rect 10320 17790 10330 17950
rect 10270 17770 10330 17790
rect 10380 17950 10440 17970
rect 10380 17790 10390 17950
rect 10430 17790 10440 17950
rect 10380 17710 10440 17790
rect 10660 17790 10670 18150
rect 10710 17790 10720 18150
rect 10660 17710 10720 17790
rect 10920 18150 10980 18310
rect 10920 17790 10930 18150
rect 10970 17790 10980 18150
rect 10920 17770 10980 17790
rect 11150 17950 11210 17970
rect 11150 17790 11160 17950
rect 11200 17790 11210 17950
rect 11150 17710 11210 17790
rect 11260 17950 11320 18310
rect 11560 18290 11620 18310
rect 11820 18250 11880 18270
rect 11820 18210 11830 18250
rect 11870 18210 11880 18250
rect 11820 18190 11880 18210
rect 11660 18150 11720 18170
rect 11260 17790 11270 17950
rect 11310 17790 11320 17950
rect 11260 17770 11320 17790
rect 11370 17950 11430 17970
rect 11370 17790 11380 17950
rect 11420 17790 11430 17950
rect 11370 17710 11430 17790
rect 11660 17790 11670 18150
rect 11710 17790 11720 18150
rect 11660 17710 11720 17790
rect 11920 18150 11980 18310
rect 11920 17790 11930 18150
rect 11970 17790 11980 18150
rect 11920 17770 11980 17790
rect 12150 17950 12210 17970
rect 12150 17790 12160 17950
rect 12200 17790 12210 17950
rect 12150 17710 12210 17790
rect 12260 17950 12320 18310
rect 12640 18290 12950 18310
rect 12990 18350 13050 19430
rect 13110 19890 13170 19910
rect 13110 19430 13120 19890
rect 13160 19430 13170 19890
rect 13110 19410 13170 19430
rect 13220 19890 13280 19970
rect 13220 19430 13230 19890
rect 13270 19430 13280 19890
rect 13220 19410 13280 19430
rect 13330 19890 13390 19910
rect 13330 19430 13340 19890
rect 13380 19430 13390 19890
rect 13210 19340 13290 19350
rect 13210 19300 13230 19340
rect 13270 19300 13290 19340
rect 13210 19290 13290 19300
rect 13210 18450 13290 18460
rect 13210 18410 13230 18450
rect 13270 18410 13290 18450
rect 13210 18400 13290 18410
rect 12990 18310 13000 18350
rect 13040 18310 13050 18350
rect 12260 17790 12270 17950
rect 12310 17790 12320 17950
rect 12260 17770 12320 17790
rect 12370 17950 12430 17970
rect 12370 17790 12380 17950
rect 12420 17790 12430 17950
rect 12370 17710 12430 17790
rect 12530 17950 12590 17970
rect 12530 17790 12540 17950
rect 12580 17790 12590 17950
rect 12530 17710 12590 17790
rect 12640 17950 12700 18290
rect 12880 18230 12940 18250
rect 12880 18070 12890 18230
rect 12930 18070 12940 18230
rect 12640 17790 12650 17950
rect 12690 17790 12700 17950
rect 12640 17770 12700 17790
rect 12750 17950 12810 17970
rect 12750 17790 12760 17950
rect 12800 17790 12810 17950
rect 12750 17710 12810 17790
rect 12880 17710 12940 18070
rect 12990 18230 13050 18310
rect 13120 18350 13180 18370
rect 13120 18310 13130 18350
rect 13170 18310 13180 18350
rect 13120 18290 13180 18310
rect 13330 18350 13390 19430
rect 13450 19890 13510 19910
rect 13450 19430 13460 19890
rect 13500 19430 13510 19890
rect 13450 19410 13510 19430
rect 13560 19890 13620 19970
rect 13560 19430 13570 19890
rect 13610 19430 13620 19890
rect 13560 19410 13620 19430
rect 13670 19890 13730 19910
rect 13670 19430 13680 19890
rect 13720 19430 13730 19890
rect 13670 19410 13730 19430
rect 13780 19890 13840 19970
rect 13780 19430 13790 19890
rect 13830 19430 13840 19890
rect 13780 19410 13840 19430
rect 13890 19890 13950 19910
rect 13890 19430 13900 19890
rect 13940 19430 13950 19890
rect 13550 19340 13630 19350
rect 13550 19300 13570 19340
rect 13610 19300 13630 19340
rect 13550 19290 13630 19300
rect 13770 19340 13850 19350
rect 13770 19300 13790 19340
rect 13830 19300 13850 19340
rect 13770 19290 13850 19300
rect 13550 18450 13630 18460
rect 13550 18410 13570 18450
rect 13610 18410 13630 18450
rect 13550 18400 13630 18410
rect 13770 18450 13850 18460
rect 13770 18410 13790 18450
rect 13830 18410 13850 18450
rect 13770 18400 13850 18410
rect 13330 18310 13340 18350
rect 13380 18310 13390 18350
rect 12990 18070 13000 18230
rect 13040 18070 13050 18230
rect 12990 18050 13050 18070
rect 13110 18230 13170 18250
rect 13110 18070 13120 18230
rect 13160 18070 13170 18230
rect 13110 18050 13170 18070
rect 13220 18230 13280 18250
rect 13220 18070 13230 18230
rect 13270 18070 13280 18230
rect 13220 17710 13280 18070
rect 13330 18230 13390 18310
rect 13460 18350 13520 18370
rect 13460 18310 13470 18350
rect 13510 18310 13520 18350
rect 13460 18290 13520 18310
rect 13890 18350 13950 19430
rect 14010 19890 14070 19910
rect 14010 19430 14020 19890
rect 14060 19430 14070 19890
rect 14010 19410 14070 19430
rect 14120 19890 14180 19970
rect 14120 19430 14130 19890
rect 14170 19430 14180 19890
rect 14120 19410 14180 19430
rect 14230 19890 14290 19910
rect 14230 19430 14240 19890
rect 14280 19430 14290 19890
rect 14230 19410 14290 19430
rect 14340 19890 14400 19970
rect 14340 19430 14350 19890
rect 14390 19430 14400 19890
rect 14340 19410 14400 19430
rect 14450 19890 14510 19910
rect 14450 19430 14460 19890
rect 14500 19430 14510 19890
rect 14450 19410 14510 19430
rect 14560 19890 14620 19970
rect 14560 19430 14570 19890
rect 14610 19430 14620 19890
rect 14560 19410 14620 19430
rect 14670 19890 14730 19910
rect 14670 19430 14680 19890
rect 14720 19430 14730 19890
rect 14670 19410 14730 19430
rect 14780 19890 14840 19970
rect 14780 19430 14790 19890
rect 14830 19430 14840 19890
rect 14780 19410 14840 19430
rect 14890 19890 14950 19910
rect 14890 19430 14900 19890
rect 14940 19430 14950 19890
rect 14110 19360 14190 19370
rect 14110 19320 14130 19360
rect 14170 19320 14190 19360
rect 14110 19310 14190 19320
rect 14330 19360 14410 19370
rect 14330 19320 14350 19360
rect 14390 19320 14410 19360
rect 14330 19310 14410 19320
rect 14550 19360 14630 19370
rect 14550 19320 14570 19360
rect 14610 19320 14630 19360
rect 14550 19310 14630 19320
rect 14770 19360 14850 19370
rect 14770 19320 14790 19360
rect 14830 19320 14850 19360
rect 14770 19310 14850 19320
rect 14110 18470 14190 18480
rect 14110 18430 14130 18470
rect 14170 18430 14190 18470
rect 14110 18420 14190 18430
rect 14330 18470 14410 18480
rect 14330 18430 14350 18470
rect 14390 18430 14410 18470
rect 14330 18420 14410 18430
rect 14550 18470 14630 18480
rect 14550 18430 14570 18470
rect 14610 18430 14630 18470
rect 14550 18420 14630 18430
rect 14770 18470 14850 18480
rect 14770 18430 14790 18470
rect 14830 18430 14850 18470
rect 14770 18420 14850 18430
rect 13890 18310 13900 18350
rect 13940 18310 13950 18350
rect 13330 18070 13340 18230
rect 13380 18070 13390 18230
rect 13330 18050 13390 18070
rect 13450 18230 13510 18250
rect 13450 18070 13460 18230
rect 13500 18070 13510 18230
rect 13450 18050 13510 18070
rect 13560 18230 13620 18250
rect 13560 18070 13570 18230
rect 13610 18070 13620 18230
rect 13560 17710 13620 18070
rect 13670 18230 13730 18250
rect 13670 18070 13680 18230
rect 13720 18070 13730 18230
rect 13670 18050 13730 18070
rect 13780 18230 13840 18250
rect 13780 18070 13790 18230
rect 13830 18070 13840 18230
rect 13780 17710 13840 18070
rect 13890 18230 13950 18310
rect 14020 18350 14080 18370
rect 14020 18310 14030 18350
rect 14070 18310 14080 18350
rect 14020 18290 14080 18310
rect 14890 18350 14950 19430
rect 15070 19890 15130 19910
rect 15070 19430 15080 19890
rect 15120 19430 15130 19890
rect 15070 19410 15130 19430
rect 15180 19890 15240 19970
rect 15180 19430 15190 19890
rect 15230 19430 15240 19890
rect 15180 19410 15240 19430
rect 15290 19890 15350 19910
rect 15290 19430 15300 19890
rect 15340 19430 15350 19890
rect 15290 19410 15350 19430
rect 15400 19890 15460 19970
rect 15400 19430 15410 19890
rect 15450 19430 15460 19890
rect 15400 19410 15460 19430
rect 15510 19890 15570 19910
rect 15510 19430 15520 19890
rect 15560 19430 15570 19890
rect 15510 19410 15570 19430
rect 15620 19890 15680 19970
rect 15620 19430 15630 19890
rect 15670 19430 15680 19890
rect 15620 19410 15680 19430
rect 15730 19890 15790 19910
rect 15730 19430 15740 19890
rect 15780 19430 15790 19890
rect 15730 19410 15790 19430
rect 15840 19890 15900 19970
rect 15840 19430 15850 19890
rect 15890 19430 15900 19890
rect 15840 19410 15900 19430
rect 15950 19890 16010 19910
rect 15950 19430 15960 19890
rect 16000 19430 16010 19890
rect 15950 19410 16010 19430
rect 16060 19890 16120 19970
rect 16060 19430 16070 19890
rect 16110 19430 16120 19890
rect 16060 19410 16120 19430
rect 16170 19890 16230 19910
rect 16170 19430 16180 19890
rect 16220 19430 16230 19890
rect 16170 19410 16230 19430
rect 16280 19890 16340 19970
rect 16280 19430 16290 19890
rect 16330 19430 16340 19890
rect 16280 19410 16340 19430
rect 16390 19890 16450 19910
rect 16390 19430 16400 19890
rect 16440 19430 16450 19890
rect 16390 19410 16450 19430
rect 16500 19890 16560 19970
rect 16500 19430 16510 19890
rect 16550 19430 16560 19890
rect 16500 19410 16560 19430
rect 16610 19890 16670 19910
rect 16610 19430 16620 19890
rect 16660 19430 16670 19890
rect 16610 19410 16670 19430
rect 16720 19890 16780 19970
rect 16720 19430 16730 19890
rect 16770 19430 16780 19890
rect 16720 19410 16780 19430
rect 16830 19890 16890 19910
rect 16830 19430 16840 19890
rect 16880 19430 16890 19890
rect 15170 19360 15250 19370
rect 15170 19320 15190 19360
rect 15230 19320 15250 19360
rect 15170 19310 15250 19320
rect 15390 19360 15470 19370
rect 15390 19320 15410 19360
rect 15450 19320 15470 19360
rect 15390 19310 15470 19320
rect 15610 19360 15690 19370
rect 15610 19320 15630 19360
rect 15670 19320 15690 19360
rect 15610 19310 15690 19320
rect 15830 19360 15910 19370
rect 15830 19320 15850 19360
rect 15890 19320 15910 19360
rect 15830 19310 15910 19320
rect 16050 19360 16130 19370
rect 16050 19320 16070 19360
rect 16110 19320 16130 19360
rect 16050 19310 16130 19320
rect 16270 19360 16350 19370
rect 16270 19320 16290 19360
rect 16330 19320 16350 19360
rect 16270 19310 16350 19320
rect 16490 19360 16570 19370
rect 16490 19320 16510 19360
rect 16550 19320 16570 19360
rect 16490 19310 16570 19320
rect 16710 19360 16790 19370
rect 16710 19320 16730 19360
rect 16770 19320 16790 19360
rect 16710 19310 16790 19320
rect 15170 18470 15250 18480
rect 15170 18430 15190 18470
rect 15230 18430 15250 18470
rect 15170 18420 15250 18430
rect 15390 18470 15470 18480
rect 15390 18430 15410 18470
rect 15450 18430 15470 18470
rect 15390 18420 15470 18430
rect 15610 18470 15690 18480
rect 15610 18430 15630 18470
rect 15670 18430 15690 18470
rect 15610 18420 15690 18430
rect 15830 18470 15910 18480
rect 15830 18430 15850 18470
rect 15890 18430 15910 18470
rect 15830 18420 15910 18430
rect 16050 18470 16130 18480
rect 16050 18430 16070 18470
rect 16110 18430 16130 18470
rect 16050 18420 16130 18430
rect 16270 18470 16350 18480
rect 16270 18430 16290 18470
rect 16330 18430 16350 18470
rect 16270 18420 16350 18430
rect 16490 18470 16570 18480
rect 16490 18430 16510 18470
rect 16550 18430 16570 18470
rect 16490 18420 16570 18430
rect 16710 18470 16790 18480
rect 16710 18430 16730 18470
rect 16770 18430 16790 18470
rect 16710 18420 16790 18430
rect 14890 18310 14900 18350
rect 14940 18310 14950 18350
rect 13890 18070 13900 18230
rect 13940 18070 13950 18230
rect 13890 18050 13950 18070
rect 14010 18230 14070 18250
rect 14010 18070 14020 18230
rect 14060 18070 14070 18230
rect 14010 18050 14070 18070
rect 14120 18230 14180 18250
rect 14120 18070 14130 18230
rect 14170 18070 14180 18230
rect 14120 17710 14180 18070
rect 14230 18230 14290 18250
rect 14230 18070 14240 18230
rect 14280 18070 14290 18230
rect 14230 18050 14290 18070
rect 14340 18230 14400 18250
rect 14340 18070 14350 18230
rect 14390 18070 14400 18230
rect 14340 17710 14400 18070
rect 14450 18230 14510 18250
rect 14450 18070 14460 18230
rect 14500 18070 14510 18230
rect 14450 18050 14510 18070
rect 14560 18230 14620 18250
rect 14560 18070 14570 18230
rect 14610 18070 14620 18230
rect 14560 17710 14620 18070
rect 14670 18230 14730 18250
rect 14670 18070 14680 18230
rect 14720 18070 14730 18230
rect 14670 18050 14730 18070
rect 14780 18230 14840 18250
rect 14780 18070 14790 18230
rect 14830 18070 14840 18230
rect 14780 17710 14840 18070
rect 14890 18230 14950 18310
rect 15080 18350 15140 18370
rect 15080 18310 15090 18350
rect 15130 18310 15140 18350
rect 15080 18290 15140 18310
rect 16830 18360 16890 19430
rect 17020 19890 17080 19910
rect 17020 19430 17030 19890
rect 17070 19430 17080 19890
rect 17020 19410 17080 19430
rect 17130 19890 17190 19970
rect 17130 19430 17140 19890
rect 17180 19430 17190 19890
rect 17130 19410 17190 19430
rect 17240 19890 17300 19910
rect 17240 19430 17250 19890
rect 17290 19430 17300 19890
rect 17240 19410 17300 19430
rect 17350 19890 17410 19970
rect 17350 19430 17360 19890
rect 17400 19430 17410 19890
rect 17350 19410 17410 19430
rect 17460 19890 17520 19910
rect 17460 19430 17470 19890
rect 17510 19430 17520 19890
rect 17460 19410 17520 19430
rect 17570 19890 17630 19970
rect 17570 19430 17580 19890
rect 17620 19430 17630 19890
rect 17570 19410 17630 19430
rect 17680 19890 17740 19910
rect 17680 19430 17690 19890
rect 17730 19430 17740 19890
rect 17680 19410 17740 19430
rect 17790 19890 17850 19970
rect 17790 19430 17800 19890
rect 17840 19430 17850 19890
rect 17790 19410 17850 19430
rect 17900 19890 17960 19910
rect 17900 19430 17910 19890
rect 17950 19430 17960 19890
rect 17900 19410 17960 19430
rect 18010 19890 18070 19970
rect 18010 19430 18020 19890
rect 18060 19430 18070 19890
rect 18010 19410 18070 19430
rect 18120 19890 18180 19910
rect 18120 19430 18130 19890
rect 18170 19430 18180 19890
rect 18120 19410 18180 19430
rect 18230 19890 18290 19970
rect 18230 19430 18240 19890
rect 18280 19430 18290 19890
rect 18230 19410 18290 19430
rect 18340 19890 18400 19910
rect 18340 19430 18350 19890
rect 18390 19430 18400 19890
rect 18340 19410 18400 19430
rect 18450 19890 18510 19970
rect 18450 19430 18460 19890
rect 18500 19430 18510 19890
rect 18450 19410 18510 19430
rect 18560 19890 18620 19910
rect 18560 19430 18570 19890
rect 18610 19430 18620 19890
rect 18560 19410 18620 19430
rect 18670 19890 18730 19970
rect 18670 19430 18680 19890
rect 18720 19430 18730 19890
rect 18670 19410 18730 19430
rect 18780 19890 18840 19910
rect 18780 19430 18790 19890
rect 18830 19430 18840 19890
rect 18780 19410 18840 19430
rect 18890 19890 18950 19970
rect 18890 19430 18900 19890
rect 18940 19430 18950 19890
rect 18890 19410 18950 19430
rect 19000 19890 19060 19910
rect 19000 19430 19010 19890
rect 19050 19430 19060 19890
rect 19000 19410 19060 19430
rect 19110 19890 19170 19970
rect 19110 19430 19120 19890
rect 19160 19430 19170 19890
rect 19110 19410 19170 19430
rect 19220 19890 19280 19910
rect 19220 19430 19230 19890
rect 19270 19430 19280 19890
rect 19220 19410 19280 19430
rect 19330 19890 19390 19970
rect 19330 19430 19340 19890
rect 19380 19430 19390 19890
rect 19330 19410 19390 19430
rect 19440 19890 19500 19910
rect 19440 19430 19450 19890
rect 19490 19430 19500 19890
rect 19440 19410 19500 19430
rect 19550 19890 19610 19970
rect 19550 19430 19560 19890
rect 19600 19430 19610 19890
rect 19550 19410 19610 19430
rect 19660 19890 19720 19910
rect 19660 19430 19670 19890
rect 19710 19430 19720 19890
rect 19660 19410 19720 19430
rect 19770 19890 19830 19970
rect 19770 19430 19780 19890
rect 19820 19430 19830 19890
rect 19770 19410 19830 19430
rect 19880 19890 19940 19910
rect 19880 19430 19890 19890
rect 19930 19430 19940 19890
rect 19880 19410 19940 19430
rect 19990 19890 20050 19970
rect 19990 19430 20000 19890
rect 20040 19430 20050 19890
rect 19990 19410 20050 19430
rect 20100 19890 20160 19910
rect 20100 19430 20110 19890
rect 20150 19430 20160 19890
rect 20100 19410 20160 19430
rect 20210 19890 20270 19970
rect 20210 19430 20220 19890
rect 20260 19430 20270 19890
rect 20210 19410 20270 19430
rect 20320 19890 20380 19910
rect 20320 19430 20330 19890
rect 20370 19430 20380 19890
rect 20320 19410 20380 19430
rect 20430 19890 20490 19970
rect 20430 19430 20440 19890
rect 20480 19430 20490 19890
rect 20430 19410 20490 19430
rect 20540 19890 20600 19910
rect 20540 19430 20550 19890
rect 20590 19430 20600 19890
rect 17120 19360 17200 19370
rect 17120 19320 17140 19360
rect 17180 19320 17200 19360
rect 17120 19310 17200 19320
rect 17340 19360 17420 19370
rect 17340 19320 17360 19360
rect 17400 19320 17420 19360
rect 17340 19310 17420 19320
rect 17560 19360 17640 19370
rect 17560 19320 17580 19360
rect 17620 19320 17640 19360
rect 17560 19310 17640 19320
rect 17780 19360 17860 19370
rect 17780 19320 17800 19360
rect 17840 19320 17860 19360
rect 17780 19310 17860 19320
rect 18000 19360 18080 19370
rect 18000 19320 18020 19360
rect 18060 19320 18080 19360
rect 18000 19310 18080 19320
rect 18220 19360 18300 19370
rect 18220 19320 18240 19360
rect 18280 19320 18300 19360
rect 18220 19310 18300 19320
rect 18440 19360 18520 19370
rect 18440 19320 18460 19360
rect 18500 19320 18520 19360
rect 18440 19310 18520 19320
rect 18660 19360 18740 19370
rect 18660 19320 18680 19360
rect 18720 19320 18740 19360
rect 18660 19310 18740 19320
rect 18880 19360 18960 19370
rect 18880 19320 18900 19360
rect 18940 19320 18960 19360
rect 18880 19310 18960 19320
rect 19100 19360 19180 19370
rect 19100 19320 19120 19360
rect 19160 19320 19180 19360
rect 19100 19310 19180 19320
rect 19320 19360 19400 19370
rect 19320 19320 19340 19360
rect 19380 19320 19400 19360
rect 19320 19310 19400 19320
rect 19540 19360 19620 19370
rect 19540 19320 19560 19360
rect 19600 19320 19620 19360
rect 19540 19310 19620 19320
rect 19760 19360 19840 19370
rect 19760 19320 19780 19360
rect 19820 19320 19840 19360
rect 19760 19310 19840 19320
rect 19980 19360 20060 19370
rect 19980 19320 20000 19360
rect 20040 19320 20060 19360
rect 19980 19310 20060 19320
rect 20200 19360 20280 19370
rect 20200 19320 20220 19360
rect 20260 19320 20280 19360
rect 20200 19310 20280 19320
rect 20420 19360 20500 19370
rect 20420 19320 20440 19360
rect 20480 19320 20500 19360
rect 20420 19310 20500 19320
rect 17120 18470 17200 18480
rect 17120 18430 17140 18470
rect 17180 18430 17200 18470
rect 17120 18420 17200 18430
rect 17340 18470 17420 18480
rect 17340 18430 17360 18470
rect 17400 18430 17420 18470
rect 17340 18420 17420 18430
rect 17560 18470 17640 18480
rect 17560 18430 17580 18470
rect 17620 18430 17640 18470
rect 17560 18420 17640 18430
rect 17780 18470 17860 18480
rect 17780 18430 17800 18470
rect 17840 18430 17860 18470
rect 17780 18420 17860 18430
rect 18000 18470 18080 18480
rect 18000 18430 18020 18470
rect 18060 18430 18080 18470
rect 18000 18420 18080 18430
rect 18220 18470 18300 18480
rect 18220 18430 18240 18470
rect 18280 18430 18300 18470
rect 18220 18420 18300 18430
rect 18440 18470 18520 18480
rect 18440 18430 18460 18470
rect 18500 18430 18520 18470
rect 18440 18420 18520 18430
rect 18660 18470 18740 18480
rect 18660 18430 18680 18470
rect 18720 18430 18740 18470
rect 18660 18420 18740 18430
rect 18880 18470 18960 18480
rect 18880 18430 18900 18470
rect 18940 18430 18960 18470
rect 18880 18420 18960 18430
rect 19100 18470 19180 18480
rect 19100 18430 19120 18470
rect 19160 18430 19180 18470
rect 19100 18420 19180 18430
rect 19320 18470 19400 18480
rect 19320 18430 19340 18470
rect 19380 18430 19400 18470
rect 19320 18420 19400 18430
rect 19540 18470 19620 18480
rect 19540 18430 19560 18470
rect 19600 18430 19620 18470
rect 19540 18420 19620 18430
rect 19760 18470 19840 18480
rect 19760 18430 19780 18470
rect 19820 18430 19840 18470
rect 19760 18420 19840 18430
rect 19980 18470 20060 18480
rect 19980 18430 20000 18470
rect 20040 18430 20060 18470
rect 19980 18420 20060 18430
rect 20200 18470 20280 18480
rect 20200 18430 20220 18470
rect 20260 18430 20280 18470
rect 20200 18420 20280 18430
rect 20420 18470 20500 18480
rect 20420 18430 20440 18470
rect 20480 18430 20500 18470
rect 20420 18420 20500 18430
rect 16830 18350 16960 18360
rect 16830 18300 16890 18350
rect 16940 18300 16960 18350
rect 16830 18290 16960 18300
rect 17020 18350 17090 18370
rect 17020 18310 17040 18350
rect 17080 18310 17090 18350
rect 17020 18290 17090 18310
rect 20540 18360 20600 19430
rect 20540 18350 20670 18360
rect 20540 18300 20600 18350
rect 20650 18300 20670 18350
rect 20540 18290 20670 18300
rect 14890 18070 14900 18230
rect 14940 18070 14950 18230
rect 14890 18050 14950 18070
rect 15070 18230 15130 18250
rect 15070 18070 15080 18230
rect 15120 18070 15130 18230
rect 15070 18050 15130 18070
rect 15180 18230 15240 18250
rect 15180 18070 15190 18230
rect 15230 18070 15240 18230
rect 15180 17710 15240 18070
rect 15290 18230 15350 18250
rect 15290 18070 15300 18230
rect 15340 18070 15350 18230
rect 15290 18050 15350 18070
rect 15400 18230 15460 18250
rect 15400 18070 15410 18230
rect 15450 18070 15460 18230
rect 15400 17710 15460 18070
rect 15510 18230 15570 18250
rect 15510 18070 15520 18230
rect 15560 18070 15570 18230
rect 15510 18050 15570 18070
rect 15620 18230 15680 18250
rect 15620 18070 15630 18230
rect 15670 18070 15680 18230
rect 15620 17710 15680 18070
rect 15730 18230 15790 18250
rect 15730 18070 15740 18230
rect 15780 18070 15790 18230
rect 15730 18050 15790 18070
rect 15840 18230 15900 18250
rect 15840 18070 15850 18230
rect 15890 18070 15900 18230
rect 15840 17710 15900 18070
rect 15950 18230 16010 18250
rect 15950 18070 15960 18230
rect 16000 18070 16010 18230
rect 15950 18050 16010 18070
rect 16060 18230 16120 18250
rect 16060 18070 16070 18230
rect 16110 18070 16120 18230
rect 16060 17710 16120 18070
rect 16170 18230 16230 18250
rect 16170 18070 16180 18230
rect 16220 18070 16230 18230
rect 16170 18050 16230 18070
rect 16280 18230 16340 18250
rect 16280 18070 16290 18230
rect 16330 18070 16340 18230
rect 16280 17710 16340 18070
rect 16390 18230 16450 18250
rect 16390 18070 16400 18230
rect 16440 18070 16450 18230
rect 16390 18050 16450 18070
rect 16500 18230 16560 18250
rect 16500 18070 16510 18230
rect 16550 18070 16560 18230
rect 16500 17710 16560 18070
rect 16610 18230 16670 18250
rect 16610 18070 16620 18230
rect 16660 18070 16670 18230
rect 16610 18050 16670 18070
rect 16720 18230 16780 18250
rect 16720 18070 16730 18230
rect 16770 18070 16780 18230
rect 16720 17710 16780 18070
rect 16830 18230 16890 18290
rect 16830 18070 16840 18230
rect 16880 18070 16890 18230
rect 16830 18050 16890 18070
rect 17020 18230 17080 18250
rect 17020 18070 17030 18230
rect 17070 18070 17080 18230
rect 17020 18050 17080 18070
rect 17130 18230 17190 18250
rect 17130 18070 17140 18230
rect 17180 18070 17190 18230
rect 17130 17710 17190 18070
rect 17240 18230 17300 18250
rect 17240 18070 17250 18230
rect 17290 18070 17300 18230
rect 17240 18050 17300 18070
rect 17350 18230 17410 18250
rect 17350 18070 17360 18230
rect 17400 18070 17410 18230
rect 17350 17710 17410 18070
rect 17460 18230 17520 18250
rect 17460 18070 17470 18230
rect 17510 18070 17520 18230
rect 17460 18050 17520 18070
rect 17570 18230 17630 18250
rect 17570 18070 17580 18230
rect 17620 18070 17630 18230
rect 17570 17710 17630 18070
rect 17680 18230 17740 18250
rect 17680 18070 17690 18230
rect 17730 18070 17740 18230
rect 17680 18050 17740 18070
rect 17790 18230 17850 18250
rect 17790 18070 17800 18230
rect 17840 18070 17850 18230
rect 17790 17710 17850 18070
rect 17900 18230 17960 18250
rect 17900 18070 17910 18230
rect 17950 18070 17960 18230
rect 17900 18050 17960 18070
rect 18010 18230 18070 18250
rect 18010 18070 18020 18230
rect 18060 18070 18070 18230
rect 18010 17710 18070 18070
rect 18120 18230 18180 18250
rect 18120 18070 18130 18230
rect 18170 18070 18180 18230
rect 18120 18050 18180 18070
rect 18230 18230 18290 18250
rect 18230 18070 18240 18230
rect 18280 18070 18290 18230
rect 18230 17710 18290 18070
rect 18340 18230 18400 18250
rect 18340 18070 18350 18230
rect 18390 18070 18400 18230
rect 18340 18050 18400 18070
rect 18450 18230 18510 18250
rect 18450 18070 18460 18230
rect 18500 18070 18510 18230
rect 18450 17710 18510 18070
rect 18560 18230 18620 18250
rect 18560 18070 18570 18230
rect 18610 18070 18620 18230
rect 18560 18050 18620 18070
rect 18670 18230 18730 18250
rect 18670 18070 18680 18230
rect 18720 18070 18730 18230
rect 18670 17710 18730 18070
rect 18780 18230 18840 18250
rect 18780 18070 18790 18230
rect 18830 18070 18840 18230
rect 18780 18050 18840 18070
rect 18890 18230 18950 18250
rect 18890 18070 18900 18230
rect 18940 18070 18950 18230
rect 18890 17710 18950 18070
rect 19000 18230 19060 18250
rect 19000 18070 19010 18230
rect 19050 18070 19060 18230
rect 19000 18050 19060 18070
rect 19110 18230 19170 18250
rect 19110 18070 19120 18230
rect 19160 18070 19170 18230
rect 19110 17710 19170 18070
rect 19220 18230 19280 18250
rect 19220 18070 19230 18230
rect 19270 18070 19280 18230
rect 19220 18050 19280 18070
rect 19330 18230 19390 18250
rect 19330 18070 19340 18230
rect 19380 18070 19390 18230
rect 19330 17710 19390 18070
rect 19440 18230 19500 18250
rect 19440 18070 19450 18230
rect 19490 18070 19500 18230
rect 19440 18050 19500 18070
rect 19550 18230 19610 18250
rect 19550 18070 19560 18230
rect 19600 18070 19610 18230
rect 19550 17710 19610 18070
rect 19660 18230 19720 18250
rect 19660 18070 19670 18230
rect 19710 18070 19720 18230
rect 19660 18050 19720 18070
rect 19770 18230 19830 18250
rect 19770 18070 19780 18230
rect 19820 18070 19830 18230
rect 19770 17710 19830 18070
rect 19880 18230 19940 18250
rect 19880 18070 19890 18230
rect 19930 18070 19940 18230
rect 19880 18050 19940 18070
rect 19990 18230 20050 18250
rect 19990 18070 20000 18230
rect 20040 18070 20050 18230
rect 19990 17710 20050 18070
rect 20100 18230 20160 18250
rect 20100 18070 20110 18230
rect 20150 18070 20160 18230
rect 20100 18050 20160 18070
rect 20210 18230 20270 18250
rect 20210 18070 20220 18230
rect 20260 18070 20270 18230
rect 20210 17710 20270 18070
rect 20320 18230 20380 18250
rect 20320 18070 20330 18230
rect 20370 18070 20380 18230
rect 20320 18050 20380 18070
rect 20430 18230 20490 18250
rect 20430 18070 20440 18230
rect 20480 18070 20490 18230
rect 20430 17710 20490 18070
rect 20540 18230 20600 18290
rect 20540 18070 20550 18230
rect 20590 18070 20600 18230
rect 20540 18050 20600 18070
rect 7280 17700 20620 17710
rect 7280 17660 7320 17700
rect 7360 17660 7400 17700
rect 7440 17660 7480 17700
rect 7520 17660 7560 17700
rect 7600 17660 7640 17700
rect 7680 17660 7720 17700
rect 7760 17660 7800 17700
rect 7840 17660 7880 17700
rect 7920 17660 7960 17700
rect 8000 17660 8040 17700
rect 8080 17660 8120 17700
rect 8160 17660 8200 17700
rect 8240 17660 8280 17700
rect 8320 17660 8360 17700
rect 8400 17660 8440 17700
rect 8480 17660 8520 17700
rect 8560 17660 8600 17700
rect 8640 17660 8680 17700
rect 8720 17660 8760 17700
rect 8800 17660 8840 17700
rect 8880 17660 8920 17700
rect 8960 17660 9000 17700
rect 9040 17660 9080 17700
rect 9120 17660 9160 17700
rect 9200 17660 9270 17700
rect 9310 17660 9350 17700
rect 9390 17660 9430 17700
rect 9470 17660 9510 17700
rect 9550 17660 9590 17700
rect 9630 17660 9670 17700
rect 9710 17660 9750 17700
rect 9790 17660 9830 17700
rect 9870 17660 9910 17700
rect 9950 17660 9990 17700
rect 10030 17660 10070 17700
rect 10110 17660 10150 17700
rect 10190 17660 10230 17700
rect 10270 17660 10310 17700
rect 10350 17660 10390 17700
rect 10430 17660 10470 17700
rect 10510 17660 10550 17700
rect 10590 17660 10630 17700
rect 10670 17660 10710 17700
rect 10750 17660 10790 17700
rect 10830 17660 10870 17700
rect 10910 17660 10950 17700
rect 10990 17660 11030 17700
rect 11070 17660 11110 17700
rect 11150 17660 11190 17700
rect 11230 17660 11270 17700
rect 11310 17660 11350 17700
rect 11390 17660 11430 17700
rect 11470 17660 11510 17700
rect 11550 17660 11590 17700
rect 11630 17660 11670 17700
rect 11710 17660 11750 17700
rect 11790 17660 11830 17700
rect 11870 17660 11910 17700
rect 11950 17660 11990 17700
rect 12030 17660 12070 17700
rect 12110 17660 12150 17700
rect 12190 17660 12230 17700
rect 12270 17660 12310 17700
rect 12350 17660 12390 17700
rect 12430 17660 12470 17700
rect 12510 17660 12550 17700
rect 12590 17660 12630 17700
rect 12670 17660 12710 17700
rect 12750 17660 12790 17700
rect 12830 17660 12870 17700
rect 12910 17660 12950 17700
rect 12990 17660 13030 17700
rect 13070 17660 13110 17700
rect 13150 17660 13190 17700
rect 13230 17660 13270 17700
rect 13310 17660 13350 17700
rect 13390 17660 13430 17700
rect 13470 17660 13510 17700
rect 13550 17660 13590 17700
rect 13630 17660 13670 17700
rect 13710 17660 13750 17700
rect 13790 17660 13830 17700
rect 13870 17660 13910 17700
rect 13950 17660 13990 17700
rect 14030 17660 14070 17700
rect 14110 17660 14150 17700
rect 14190 17660 14230 17700
rect 14270 17660 14310 17700
rect 14350 17660 14390 17700
rect 14430 17660 14470 17700
rect 14510 17660 14550 17700
rect 14590 17660 14630 17700
rect 14670 17660 14710 17700
rect 14750 17660 14790 17700
rect 14830 17660 14870 17700
rect 14910 17660 14950 17700
rect 14990 17660 15030 17700
rect 15070 17660 15110 17700
rect 15150 17660 15190 17700
rect 15230 17660 15270 17700
rect 15310 17660 15350 17700
rect 15390 17660 15430 17700
rect 15470 17660 15510 17700
rect 15550 17660 15590 17700
rect 15630 17660 15670 17700
rect 15710 17660 15750 17700
rect 15790 17660 15830 17700
rect 15870 17660 15910 17700
rect 15950 17660 15990 17700
rect 16030 17660 16070 17700
rect 16110 17660 16150 17700
rect 16190 17660 16230 17700
rect 16270 17660 16310 17700
rect 16350 17660 16390 17700
rect 16430 17660 16470 17700
rect 16510 17660 16550 17700
rect 16590 17660 16630 17700
rect 16670 17660 16710 17700
rect 16750 17660 16790 17700
rect 16830 17660 16870 17700
rect 16910 17660 16950 17700
rect 16990 17660 17030 17700
rect 17070 17660 17110 17700
rect 17150 17660 17190 17700
rect 17230 17660 17270 17700
rect 17310 17660 17350 17700
rect 17390 17660 17430 17700
rect 17470 17660 17510 17700
rect 17550 17660 17590 17700
rect 17630 17660 17670 17700
rect 17710 17660 17750 17700
rect 17790 17660 17830 17700
rect 17870 17660 17910 17700
rect 17950 17660 17990 17700
rect 18030 17660 18070 17700
rect 18110 17660 18150 17700
rect 18190 17660 18230 17700
rect 18270 17660 18310 17700
rect 18350 17660 18390 17700
rect 18430 17660 18470 17700
rect 18510 17660 18550 17700
rect 18590 17660 18630 17700
rect 18670 17660 18710 17700
rect 18750 17660 18790 17700
rect 18830 17660 18870 17700
rect 18910 17660 18950 17700
rect 18990 17660 19030 17700
rect 19070 17660 19110 17700
rect 19150 17660 19190 17700
rect 19230 17660 19270 17700
rect 19310 17660 19350 17700
rect 19390 17660 19430 17700
rect 19470 17660 19510 17700
rect 19550 17660 19590 17700
rect 19630 17660 19670 17700
rect 19710 17660 19750 17700
rect 19790 17660 19830 17700
rect 19870 17660 19910 17700
rect 19950 17660 19990 17700
rect 20030 17660 20070 17700
rect 20110 17660 20150 17700
rect 20190 17660 20230 17700
rect 20270 17660 20310 17700
rect 20350 17660 20390 17700
rect 20430 17660 20470 17700
rect 20510 17660 20550 17700
rect 20590 17660 20620 17700
rect 7280 17650 20620 17660
rect 9620 15660 21160 15670
rect 9620 15620 9710 15660
rect 9750 15620 9790 15660
rect 9830 15620 9870 15660
rect 9910 15620 9950 15660
rect 9990 15620 10030 15660
rect 10070 15620 10110 15660
rect 10150 15620 10190 15660
rect 10230 15620 10270 15660
rect 10310 15620 10350 15660
rect 10390 15620 10430 15660
rect 10470 15620 10510 15660
rect 10550 15620 10590 15660
rect 10630 15620 10670 15660
rect 10710 15620 10750 15660
rect 10790 15620 10830 15660
rect 10870 15620 10910 15660
rect 10950 15620 10990 15660
rect 11030 15620 11070 15660
rect 11110 15620 11150 15660
rect 11190 15620 11230 15660
rect 11270 15620 11310 15660
rect 11350 15620 11390 15660
rect 11430 15620 11470 15660
rect 11510 15620 11550 15660
rect 11590 15620 11630 15660
rect 11670 15620 11710 15660
rect 11750 15620 11790 15660
rect 11830 15620 11870 15660
rect 11910 15620 11950 15660
rect 11990 15620 12030 15660
rect 12070 15620 12110 15660
rect 12150 15620 12190 15660
rect 12230 15620 12270 15660
rect 12310 15620 12350 15660
rect 12390 15620 12430 15660
rect 12470 15620 12510 15660
rect 12550 15620 12590 15660
rect 12630 15620 12670 15660
rect 12710 15620 12750 15660
rect 12790 15620 12830 15660
rect 12870 15620 12910 15660
rect 12950 15620 12990 15660
rect 13030 15620 13070 15660
rect 13110 15620 13150 15660
rect 13190 15620 13230 15660
rect 13270 15620 13310 15660
rect 13350 15620 13390 15660
rect 13430 15620 13470 15660
rect 13510 15620 13550 15660
rect 13590 15620 13630 15660
rect 13670 15620 13710 15660
rect 13750 15620 13790 15660
rect 13830 15620 13870 15660
rect 13910 15620 13950 15660
rect 13990 15620 14030 15660
rect 14070 15620 14110 15660
rect 14150 15620 14190 15660
rect 14230 15620 14270 15660
rect 14310 15620 14350 15660
rect 14390 15620 14430 15660
rect 14470 15620 14510 15660
rect 14550 15620 14590 15660
rect 14630 15620 14670 15660
rect 14710 15620 14750 15660
rect 14790 15620 14830 15660
rect 14870 15620 14910 15660
rect 14950 15620 14990 15660
rect 15030 15620 15070 15660
rect 15110 15620 15150 15660
rect 15190 15620 15230 15660
rect 15270 15620 15310 15660
rect 15350 15620 15390 15660
rect 15430 15620 15470 15660
rect 15510 15620 15550 15660
rect 15590 15620 15630 15660
rect 15670 15620 15710 15660
rect 15750 15620 15790 15660
rect 15830 15620 15870 15660
rect 15910 15620 15950 15660
rect 15990 15620 16030 15660
rect 16070 15620 16110 15660
rect 16150 15620 16190 15660
rect 16230 15620 16270 15660
rect 16310 15620 16350 15660
rect 16390 15620 16430 15660
rect 16470 15620 16510 15660
rect 16550 15620 16590 15660
rect 16630 15620 16670 15660
rect 16710 15620 16750 15660
rect 16790 15620 16830 15660
rect 16870 15620 16910 15660
rect 16950 15620 16990 15660
rect 17030 15620 17070 15660
rect 17110 15620 17150 15660
rect 17190 15620 17230 15660
rect 17270 15620 17310 15660
rect 17350 15620 17390 15660
rect 17430 15620 17470 15660
rect 17510 15620 17550 15660
rect 17590 15620 17630 15660
rect 17670 15620 17710 15660
rect 17750 15620 17790 15660
rect 17830 15620 17870 15660
rect 17910 15620 17950 15660
rect 17990 15620 18030 15660
rect 18070 15620 18110 15660
rect 18150 15620 18190 15660
rect 18230 15620 18270 15660
rect 18310 15620 18350 15660
rect 18390 15620 18430 15660
rect 18470 15620 18510 15660
rect 18550 15620 18590 15660
rect 18630 15620 18670 15660
rect 18710 15620 18750 15660
rect 18790 15620 18830 15660
rect 18870 15620 18910 15660
rect 18950 15620 18990 15660
rect 19030 15620 19070 15660
rect 19110 15620 19150 15660
rect 19190 15620 19230 15660
rect 19270 15620 19310 15660
rect 19350 15620 19390 15660
rect 19430 15620 19470 15660
rect 19510 15620 19550 15660
rect 19590 15620 19630 15660
rect 19670 15620 19710 15660
rect 19750 15620 19800 15660
rect 19840 15620 19880 15660
rect 19920 15620 19960 15660
rect 20000 15620 20040 15660
rect 20080 15620 20120 15660
rect 20160 15620 20200 15660
rect 20240 15620 20280 15660
rect 20320 15620 20370 15660
rect 20410 15620 20450 15660
rect 20490 15620 20530 15660
rect 20570 15620 20610 15660
rect 20650 15620 20690 15660
rect 20730 15620 20770 15660
rect 20810 15620 20850 15660
rect 20890 15620 20930 15660
rect 20970 15620 21010 15660
rect 21050 15620 21090 15660
rect 21130 15620 21160 15660
rect 9620 15610 21160 15620
rect 9760 15530 9820 15610
rect 9760 15370 9770 15530
rect 9810 15370 9820 15530
rect 9760 15350 9820 15370
rect 9870 15530 9930 15550
rect 9870 15370 9880 15530
rect 9920 15370 9930 15530
rect 9730 15110 9830 15120
rect 9730 15050 9750 15110
rect 9810 15050 9830 15110
rect 9730 15040 9830 15050
rect 9870 15010 9930 15370
rect 9980 15530 10040 15610
rect 9980 15370 9990 15530
rect 10030 15370 10040 15530
rect 9980 15350 10040 15370
rect 10410 15530 10470 15610
rect 10410 15170 10420 15530
rect 10460 15170 10470 15530
rect 10410 15150 10470 15170
rect 10670 15530 10730 15550
rect 10670 15170 10680 15530
rect 10720 15170 10730 15530
rect 10900 15530 10960 15610
rect 10900 15370 10910 15530
rect 10950 15370 10960 15530
rect 10900 15350 10960 15370
rect 11010 15530 11070 15550
rect 11010 15370 11020 15530
rect 11060 15370 11070 15530
rect 10570 15110 10630 15130
rect 10570 15070 10580 15110
rect 10620 15070 10630 15110
rect 10570 15050 10630 15070
rect 10260 15020 10370 15030
rect 9870 15000 10120 15010
rect 9870 14960 10060 15000
rect 10100 14960 10120 15000
rect 9870 14950 10120 14960
rect 10260 14960 10280 15020
rect 10350 14960 10370 15020
rect 10670 15010 10730 15170
rect 11010 15010 11070 15370
rect 11120 15530 11180 15610
rect 11120 15370 11130 15530
rect 11170 15370 11180 15530
rect 11120 15350 11180 15370
rect 11400 15530 11460 15610
rect 11400 15170 11410 15530
rect 11450 15170 11460 15530
rect 11400 15150 11460 15170
rect 11660 15530 11720 15550
rect 11660 15170 11670 15530
rect 11710 15170 11720 15530
rect 11890 15530 11950 15610
rect 11890 15370 11900 15530
rect 11940 15370 11950 15530
rect 11890 15350 11950 15370
rect 12000 15530 12060 15550
rect 12000 15370 12010 15530
rect 12050 15370 12060 15530
rect 11560 15110 11620 15130
rect 11560 15070 11570 15110
rect 11610 15070 11620 15110
rect 11560 15050 11620 15070
rect 11300 15010 11360 15030
rect 11660 15010 11720 15170
rect 12000 15010 12060 15370
rect 12110 15530 12170 15610
rect 12110 15370 12120 15530
rect 12160 15370 12170 15530
rect 12110 15350 12170 15370
rect 12400 15530 12460 15610
rect 12400 15170 12410 15530
rect 12450 15170 12460 15530
rect 12400 15150 12460 15170
rect 12660 15530 12720 15550
rect 12660 15170 12670 15530
rect 12710 15170 12720 15530
rect 12890 15530 12950 15610
rect 12890 15370 12900 15530
rect 12940 15370 12950 15530
rect 12890 15350 12950 15370
rect 13000 15530 13060 15550
rect 13000 15370 13010 15530
rect 13050 15370 13060 15530
rect 12560 15110 12620 15130
rect 12560 15070 12570 15110
rect 12610 15070 12620 15110
rect 12560 15050 12620 15070
rect 12300 15010 12360 15030
rect 12660 15010 12720 15170
rect 13000 15030 13060 15370
rect 13110 15530 13170 15610
rect 13110 15370 13120 15530
rect 13160 15370 13170 15530
rect 13110 15350 13170 15370
rect 13240 15250 13300 15610
rect 13240 15090 13250 15250
rect 13290 15090 13300 15250
rect 13240 15070 13300 15090
rect 13350 15250 13410 15270
rect 13350 15090 13360 15250
rect 13400 15090 13410 15250
rect 13000 15010 13310 15030
rect 10260 14950 10370 14960
rect 10540 15000 10970 15010
rect 10540 14960 10820 15000
rect 10860 14960 10900 15000
rect 10940 14960 10970 15000
rect 10540 14950 10970 14960
rect 11010 15000 11250 15010
rect 11010 14960 11200 15000
rect 11240 14960 11250 15000
rect 11010 14950 11250 14960
rect 11300 14970 11310 15010
rect 11350 14970 11360 15010
rect 11300 14950 11360 14970
rect 11530 15000 11960 15010
rect 11530 14960 11810 15000
rect 11850 14960 11890 15000
rect 11930 14960 11960 15000
rect 11530 14950 11960 14960
rect 12000 15000 12240 15010
rect 12000 14960 12190 15000
rect 12230 14960 12240 15000
rect 12000 14950 12240 14960
rect 12300 14970 12310 15010
rect 12350 14970 12360 15010
rect 12300 14950 12360 14970
rect 12530 15000 12960 15010
rect 12530 14960 12810 15000
rect 12850 14960 12890 15000
rect 12930 14960 12960 15000
rect 12530 14950 12960 14960
rect 13000 14970 13180 15010
rect 13220 14970 13260 15010
rect 13300 14970 13310 15010
rect 13000 14950 13310 14970
rect 13350 15010 13410 15090
rect 13470 15250 13530 15270
rect 13470 15090 13480 15250
rect 13520 15090 13530 15250
rect 13470 15070 13530 15090
rect 13580 15250 13640 15610
rect 13580 15090 13590 15250
rect 13630 15090 13640 15250
rect 13580 15070 13640 15090
rect 13690 15250 13750 15270
rect 13690 15090 13700 15250
rect 13740 15090 13750 15250
rect 13350 14970 13360 15010
rect 13400 14970 13410 15010
rect 9760 14890 9820 14910
rect 9760 14430 9770 14890
rect 9810 14430 9820 14890
rect 9760 14350 9820 14430
rect 9870 14890 9930 14950
rect 9870 14430 9880 14890
rect 9920 14430 9930 14890
rect 9870 14410 9930 14430
rect 9980 14890 10040 14910
rect 9980 14430 9990 14890
rect 10030 14430 10040 14890
rect 9980 14350 10040 14430
rect 10410 14890 10470 14910
rect 10410 14430 10420 14890
rect 10460 14430 10470 14890
rect 10410 14350 10470 14430
rect 10540 14890 10600 14950
rect 10540 14430 10550 14890
rect 10590 14430 10600 14890
rect 10540 14410 10600 14430
rect 10670 14890 10730 14910
rect 10670 14430 10680 14890
rect 10720 14430 10730 14890
rect 10670 14350 10730 14430
rect 10900 14890 10960 14910
rect 10900 14430 10910 14890
rect 10950 14430 10960 14890
rect 10900 14350 10960 14430
rect 11010 14890 11070 14950
rect 11010 14430 11020 14890
rect 11060 14430 11070 14890
rect 11010 14410 11070 14430
rect 11120 14890 11180 14910
rect 11120 14430 11130 14890
rect 11170 14430 11180 14890
rect 11120 14350 11180 14430
rect 11400 14890 11460 14910
rect 11400 14430 11410 14890
rect 11450 14430 11460 14890
rect 11400 14350 11460 14430
rect 11530 14890 11590 14950
rect 11530 14430 11540 14890
rect 11580 14430 11590 14890
rect 11530 14410 11590 14430
rect 11660 14890 11720 14910
rect 11660 14430 11670 14890
rect 11710 14430 11720 14890
rect 11660 14350 11720 14430
rect 11890 14890 11950 14910
rect 11890 14430 11900 14890
rect 11940 14430 11950 14890
rect 11890 14350 11950 14430
rect 12000 14890 12060 14950
rect 12000 14430 12010 14890
rect 12050 14430 12060 14890
rect 12000 14410 12060 14430
rect 12110 14890 12170 14910
rect 12110 14430 12120 14890
rect 12160 14430 12170 14890
rect 12110 14350 12170 14430
rect 12400 14890 12460 14910
rect 12400 14430 12410 14890
rect 12450 14430 12460 14890
rect 12400 14350 12460 14430
rect 12530 14890 12590 14950
rect 12530 14430 12540 14890
rect 12580 14430 12590 14890
rect 12530 14410 12590 14430
rect 12660 14890 12720 14910
rect 12660 14430 12670 14890
rect 12710 14430 12720 14890
rect 12660 14350 12720 14430
rect 12890 14890 12950 14910
rect 12890 14430 12900 14890
rect 12940 14430 12950 14890
rect 12890 14350 12950 14430
rect 13000 14890 13060 14950
rect 13000 14430 13010 14890
rect 13050 14430 13060 14890
rect 13000 14410 13060 14430
rect 13110 14890 13170 14910
rect 13110 14430 13120 14890
rect 13160 14430 13170 14890
rect 13110 14350 13170 14430
rect 13240 14890 13300 14910
rect 13240 14430 13250 14890
rect 13290 14430 13300 14890
rect 13240 14350 13300 14430
rect 13350 14890 13410 14970
rect 13480 15010 13540 15030
rect 13480 14970 13490 15010
rect 13530 14970 13540 15010
rect 13480 14950 13540 14970
rect 13690 15010 13750 15090
rect 13810 15250 13870 15270
rect 13810 15090 13820 15250
rect 13860 15090 13870 15250
rect 13810 15070 13870 15090
rect 13920 15250 13980 15610
rect 13920 15090 13930 15250
rect 13970 15090 13980 15250
rect 13920 15070 13980 15090
rect 14030 15250 14090 15270
rect 14030 15090 14040 15250
rect 14080 15090 14090 15250
rect 14030 15070 14090 15090
rect 14140 15250 14200 15610
rect 14140 15090 14150 15250
rect 14190 15090 14200 15250
rect 14140 15070 14200 15090
rect 14250 15250 14310 15270
rect 14250 15090 14260 15250
rect 14300 15090 14310 15250
rect 13690 14970 13700 15010
rect 13740 14970 13750 15010
rect 13350 14430 13360 14890
rect 13400 14430 13410 14890
rect 13350 14410 13410 14430
rect 13470 14890 13530 14910
rect 13470 14430 13480 14890
rect 13520 14430 13530 14890
rect 13470 14410 13530 14430
rect 13580 14890 13640 14910
rect 13580 14430 13590 14890
rect 13630 14430 13640 14890
rect 13580 14350 13640 14430
rect 13690 14890 13750 14970
rect 13820 15010 13880 15030
rect 13820 14970 13830 15010
rect 13870 14970 13880 15010
rect 13820 14950 13880 14970
rect 14250 15010 14310 15090
rect 14370 15250 14430 15270
rect 14370 15090 14380 15250
rect 14420 15090 14430 15250
rect 14370 15070 14430 15090
rect 14480 15250 14540 15610
rect 14480 15090 14490 15250
rect 14530 15090 14540 15250
rect 14480 15070 14540 15090
rect 14590 15250 14650 15270
rect 14590 15090 14600 15250
rect 14640 15090 14650 15250
rect 14590 15070 14650 15090
rect 14700 15250 14760 15610
rect 14700 15090 14710 15250
rect 14750 15090 14760 15250
rect 14700 15070 14760 15090
rect 14810 15250 14870 15270
rect 14810 15090 14820 15250
rect 14860 15090 14870 15250
rect 14810 15070 14870 15090
rect 14920 15250 14980 15610
rect 14920 15090 14930 15250
rect 14970 15090 14980 15250
rect 14920 15070 14980 15090
rect 15030 15250 15090 15270
rect 15030 15090 15040 15250
rect 15080 15090 15090 15250
rect 15030 15070 15090 15090
rect 15140 15250 15200 15610
rect 15140 15090 15150 15250
rect 15190 15090 15200 15250
rect 15140 15070 15200 15090
rect 15250 15250 15310 15270
rect 15250 15090 15260 15250
rect 15300 15090 15310 15250
rect 14250 14970 14260 15010
rect 14300 14970 14310 15010
rect 13690 14430 13700 14890
rect 13740 14430 13750 14890
rect 13690 14410 13750 14430
rect 13810 14890 13870 14910
rect 13810 14430 13820 14890
rect 13860 14430 13870 14890
rect 13810 14410 13870 14430
rect 13920 14890 13980 14910
rect 13920 14430 13930 14890
rect 13970 14430 13980 14890
rect 13920 14350 13980 14430
rect 14030 14890 14090 14910
rect 14030 14430 14040 14890
rect 14080 14430 14090 14890
rect 14030 14410 14090 14430
rect 14140 14890 14200 14910
rect 14140 14430 14150 14890
rect 14190 14430 14200 14890
rect 14140 14350 14200 14430
rect 14250 14890 14310 14970
rect 14380 15010 14440 15030
rect 14380 14970 14390 15010
rect 14430 14970 14440 15010
rect 14380 14950 14440 14970
rect 15250 15010 15310 15090
rect 15430 15250 15490 15270
rect 15430 15090 15440 15250
rect 15480 15090 15490 15250
rect 15430 15070 15490 15090
rect 15540 15250 15600 15610
rect 15540 15090 15550 15250
rect 15590 15090 15600 15250
rect 15540 15070 15600 15090
rect 15650 15250 15710 15270
rect 15650 15090 15660 15250
rect 15700 15090 15710 15250
rect 15650 15070 15710 15090
rect 15760 15250 15820 15610
rect 15760 15090 15770 15250
rect 15810 15090 15820 15250
rect 15760 15070 15820 15090
rect 15870 15250 15930 15270
rect 15870 15090 15880 15250
rect 15920 15090 15930 15250
rect 15870 15070 15930 15090
rect 15980 15250 16040 15610
rect 15980 15090 15990 15250
rect 16030 15090 16040 15250
rect 15980 15070 16040 15090
rect 16090 15250 16150 15270
rect 16090 15090 16100 15250
rect 16140 15090 16150 15250
rect 16090 15070 16150 15090
rect 16200 15250 16260 15610
rect 16200 15090 16210 15250
rect 16250 15090 16260 15250
rect 16200 15070 16260 15090
rect 16310 15250 16370 15270
rect 16310 15090 16320 15250
rect 16360 15090 16370 15250
rect 16310 15070 16370 15090
rect 16420 15250 16480 15610
rect 16420 15090 16430 15250
rect 16470 15090 16480 15250
rect 16420 15070 16480 15090
rect 16530 15250 16590 15270
rect 16530 15090 16540 15250
rect 16580 15090 16590 15250
rect 16530 15070 16590 15090
rect 16640 15250 16700 15610
rect 16640 15090 16650 15250
rect 16690 15090 16700 15250
rect 16640 15070 16700 15090
rect 16750 15250 16810 15270
rect 16750 15090 16760 15250
rect 16800 15090 16810 15250
rect 16750 15070 16810 15090
rect 16860 15250 16920 15610
rect 16860 15090 16870 15250
rect 16910 15090 16920 15250
rect 16860 15070 16920 15090
rect 16970 15250 17030 15270
rect 16970 15090 16980 15250
rect 17020 15090 17030 15250
rect 16970 15070 17030 15090
rect 17080 15250 17140 15610
rect 17080 15090 17090 15250
rect 17130 15090 17140 15250
rect 17080 15070 17140 15090
rect 17190 15250 17250 15270
rect 17190 15090 17200 15250
rect 17240 15090 17250 15250
rect 17190 15030 17250 15090
rect 17380 15250 17440 15270
rect 17380 15090 17390 15250
rect 17430 15090 17440 15250
rect 17380 15070 17440 15090
rect 17490 15250 17550 15610
rect 17490 15090 17500 15250
rect 17540 15090 17550 15250
rect 17490 15070 17550 15090
rect 17600 15250 17660 15270
rect 17600 15090 17610 15250
rect 17650 15090 17660 15250
rect 17600 15070 17660 15090
rect 17710 15250 17770 15610
rect 17710 15090 17720 15250
rect 17760 15090 17770 15250
rect 17710 15070 17770 15090
rect 17820 15250 17880 15270
rect 17820 15090 17830 15250
rect 17870 15090 17880 15250
rect 17820 15070 17880 15090
rect 17930 15250 17990 15610
rect 17930 15090 17940 15250
rect 17980 15090 17990 15250
rect 17930 15070 17990 15090
rect 18040 15250 18100 15270
rect 18040 15090 18050 15250
rect 18090 15090 18100 15250
rect 18040 15070 18100 15090
rect 18150 15250 18210 15610
rect 18150 15090 18160 15250
rect 18200 15090 18210 15250
rect 18150 15070 18210 15090
rect 18260 15250 18320 15270
rect 18260 15090 18270 15250
rect 18310 15090 18320 15250
rect 18260 15070 18320 15090
rect 18370 15250 18430 15610
rect 18370 15090 18380 15250
rect 18420 15090 18430 15250
rect 18370 15070 18430 15090
rect 18480 15250 18540 15270
rect 18480 15090 18490 15250
rect 18530 15090 18540 15250
rect 18480 15070 18540 15090
rect 18590 15250 18650 15610
rect 18590 15090 18600 15250
rect 18640 15090 18650 15250
rect 18590 15070 18650 15090
rect 18700 15250 18760 15270
rect 18700 15090 18710 15250
rect 18750 15090 18760 15250
rect 18700 15070 18760 15090
rect 18810 15250 18870 15610
rect 18810 15090 18820 15250
rect 18860 15090 18870 15250
rect 18810 15070 18870 15090
rect 18920 15250 18980 15270
rect 18920 15090 18930 15250
rect 18970 15090 18980 15250
rect 18920 15070 18980 15090
rect 19030 15250 19090 15610
rect 19030 15090 19040 15250
rect 19080 15090 19090 15250
rect 19030 15070 19090 15090
rect 19140 15250 19200 15270
rect 19140 15090 19150 15250
rect 19190 15090 19200 15250
rect 19140 15070 19200 15090
rect 19250 15250 19310 15610
rect 19250 15090 19260 15250
rect 19300 15090 19310 15250
rect 19250 15070 19310 15090
rect 19360 15250 19420 15270
rect 19360 15090 19370 15250
rect 19410 15090 19420 15250
rect 19360 15070 19420 15090
rect 19470 15250 19530 15610
rect 19470 15090 19480 15250
rect 19520 15090 19530 15250
rect 19470 15070 19530 15090
rect 19580 15250 19640 15270
rect 19580 15090 19590 15250
rect 19630 15090 19640 15250
rect 19580 15070 19640 15090
rect 19690 15250 19750 15610
rect 19690 15090 19700 15250
rect 19740 15090 19750 15250
rect 19690 15070 19750 15090
rect 19800 15250 19860 15270
rect 19800 15090 19810 15250
rect 19850 15090 19860 15250
rect 19800 15070 19860 15090
rect 19910 15250 19970 15610
rect 19910 15090 19920 15250
rect 19960 15090 19970 15250
rect 19910 15070 19970 15090
rect 20020 15250 20080 15270
rect 20020 15090 20030 15250
rect 20070 15090 20080 15250
rect 20020 15070 20080 15090
rect 20130 15250 20190 15610
rect 20130 15090 20140 15250
rect 20180 15090 20190 15250
rect 20130 15070 20190 15090
rect 20240 15250 20300 15270
rect 20240 15090 20250 15250
rect 20290 15090 20300 15250
rect 20240 15070 20300 15090
rect 20350 15250 20410 15610
rect 20350 15090 20360 15250
rect 20400 15090 20410 15250
rect 20350 15070 20410 15090
rect 20460 15250 20520 15270
rect 20460 15090 20470 15250
rect 20510 15090 20520 15250
rect 20460 15070 20520 15090
rect 20570 15250 20630 15610
rect 20570 15090 20580 15250
rect 20620 15090 20630 15250
rect 20570 15070 20630 15090
rect 20680 15250 20740 15270
rect 20680 15090 20690 15250
rect 20730 15090 20740 15250
rect 20680 15070 20740 15090
rect 20790 15250 20850 15610
rect 20790 15090 20800 15250
rect 20840 15090 20850 15250
rect 20790 15070 20850 15090
rect 20900 15250 20960 15270
rect 20900 15090 20910 15250
rect 20950 15090 20960 15250
rect 20900 15030 20960 15090
rect 15250 14970 15260 15010
rect 15300 14970 15310 15010
rect 14250 14430 14260 14890
rect 14300 14430 14310 14890
rect 14250 14410 14310 14430
rect 14370 14890 14430 14910
rect 14370 14430 14380 14890
rect 14420 14430 14430 14890
rect 14370 14410 14430 14430
rect 14480 14890 14540 14910
rect 14480 14430 14490 14890
rect 14530 14430 14540 14890
rect 14480 14350 14540 14430
rect 14590 14890 14650 14910
rect 14590 14430 14600 14890
rect 14640 14430 14650 14890
rect 14590 14410 14650 14430
rect 14700 14890 14760 14910
rect 14700 14430 14710 14890
rect 14750 14430 14760 14890
rect 14700 14350 14760 14430
rect 14810 14890 14870 14910
rect 14810 14430 14820 14890
rect 14860 14430 14870 14890
rect 14810 14410 14870 14430
rect 14920 14890 14980 14910
rect 14920 14430 14930 14890
rect 14970 14430 14980 14890
rect 14920 14350 14980 14430
rect 15030 14890 15090 14910
rect 15030 14430 15040 14890
rect 15080 14430 15090 14890
rect 15030 14410 15090 14430
rect 15140 14890 15200 14910
rect 15140 14430 15150 14890
rect 15190 14430 15200 14890
rect 15140 14350 15200 14430
rect 15250 14890 15310 14970
rect 15440 15010 15500 15030
rect 15440 14970 15450 15010
rect 15490 14970 15500 15010
rect 15440 14950 15500 14970
rect 17190 15020 17320 15030
rect 17190 14970 17250 15020
rect 17300 14970 17320 15020
rect 17190 14960 17320 14970
rect 17380 15010 17450 15030
rect 17380 14970 17400 15010
rect 17440 14970 17450 15010
rect 15250 14430 15260 14890
rect 15300 14430 15310 14890
rect 15250 14410 15310 14430
rect 15430 14890 15490 14910
rect 15430 14430 15440 14890
rect 15480 14430 15490 14890
rect 15430 14410 15490 14430
rect 15540 14890 15600 14910
rect 15540 14430 15550 14890
rect 15590 14430 15600 14890
rect 15540 14350 15600 14430
rect 15650 14890 15710 14910
rect 15650 14430 15660 14890
rect 15700 14430 15710 14890
rect 15650 14410 15710 14430
rect 15760 14890 15820 14910
rect 15760 14430 15770 14890
rect 15810 14430 15820 14890
rect 15760 14350 15820 14430
rect 15870 14890 15930 14910
rect 15870 14430 15880 14890
rect 15920 14430 15930 14890
rect 15870 14410 15930 14430
rect 15980 14890 16040 14910
rect 15980 14430 15990 14890
rect 16030 14430 16040 14890
rect 15980 14350 16040 14430
rect 16090 14890 16150 14910
rect 16090 14430 16100 14890
rect 16140 14430 16150 14890
rect 16090 14410 16150 14430
rect 16200 14890 16260 14910
rect 16200 14430 16210 14890
rect 16250 14430 16260 14890
rect 16200 14350 16260 14430
rect 16310 14890 16370 14910
rect 16310 14430 16320 14890
rect 16360 14430 16370 14890
rect 16310 14410 16370 14430
rect 16420 14890 16480 14910
rect 16420 14430 16430 14890
rect 16470 14430 16480 14890
rect 16420 14350 16480 14430
rect 16530 14890 16590 14910
rect 16530 14430 16540 14890
rect 16580 14430 16590 14890
rect 16530 14410 16590 14430
rect 16640 14890 16700 14910
rect 16640 14430 16650 14890
rect 16690 14430 16700 14890
rect 16640 14350 16700 14430
rect 16750 14890 16810 14910
rect 16750 14430 16760 14890
rect 16800 14430 16810 14890
rect 16750 14410 16810 14430
rect 16860 14890 16920 14910
rect 16860 14430 16870 14890
rect 16910 14430 16920 14890
rect 16860 14350 16920 14430
rect 16970 14890 17030 14910
rect 16970 14430 16980 14890
rect 17020 14430 17030 14890
rect 16970 14410 17030 14430
rect 17080 14890 17140 14910
rect 17080 14430 17090 14890
rect 17130 14430 17140 14890
rect 17080 14350 17140 14430
rect 17190 14890 17250 14960
rect 17380 14950 17450 14970
rect 20900 15020 21030 15030
rect 20900 14970 20960 15020
rect 21010 14970 21030 15020
rect 20900 14960 21030 14970
rect 17190 14430 17200 14890
rect 17240 14430 17250 14890
rect 17190 14410 17250 14430
rect 17380 14890 17440 14910
rect 17380 14430 17390 14890
rect 17430 14430 17440 14890
rect 17380 14410 17440 14430
rect 17490 14890 17550 14910
rect 17490 14430 17500 14890
rect 17540 14430 17550 14890
rect 17490 14350 17550 14430
rect 17600 14890 17660 14910
rect 17600 14430 17610 14890
rect 17650 14430 17660 14890
rect 17600 14410 17660 14430
rect 17710 14890 17770 14910
rect 17710 14430 17720 14890
rect 17760 14430 17770 14890
rect 17710 14350 17770 14430
rect 17820 14890 17880 14910
rect 17820 14430 17830 14890
rect 17870 14430 17880 14890
rect 17820 14410 17880 14430
rect 17930 14890 17990 14910
rect 17930 14430 17940 14890
rect 17980 14430 17990 14890
rect 17930 14350 17990 14430
rect 18040 14890 18100 14910
rect 18040 14430 18050 14890
rect 18090 14430 18100 14890
rect 18040 14410 18100 14430
rect 18150 14890 18210 14910
rect 18150 14430 18160 14890
rect 18200 14430 18210 14890
rect 18150 14350 18210 14430
rect 18260 14890 18320 14910
rect 18260 14430 18270 14890
rect 18310 14430 18320 14890
rect 18260 14410 18320 14430
rect 18370 14890 18430 14910
rect 18370 14430 18380 14890
rect 18420 14430 18430 14890
rect 18370 14350 18430 14430
rect 18480 14890 18540 14910
rect 18480 14430 18490 14890
rect 18530 14430 18540 14890
rect 18480 14410 18540 14430
rect 18590 14890 18650 14910
rect 18590 14430 18600 14890
rect 18640 14430 18650 14890
rect 18590 14350 18650 14430
rect 18700 14890 18760 14910
rect 18700 14430 18710 14890
rect 18750 14430 18760 14890
rect 18700 14410 18760 14430
rect 18810 14890 18870 14910
rect 18810 14430 18820 14890
rect 18860 14430 18870 14890
rect 18810 14350 18870 14430
rect 18920 14890 18980 14910
rect 18920 14430 18930 14890
rect 18970 14430 18980 14890
rect 18920 14410 18980 14430
rect 19030 14890 19090 14910
rect 19030 14430 19040 14890
rect 19080 14430 19090 14890
rect 19030 14350 19090 14430
rect 19140 14890 19200 14910
rect 19140 14430 19150 14890
rect 19190 14430 19200 14890
rect 19140 14410 19200 14430
rect 19250 14890 19310 14910
rect 19250 14430 19260 14890
rect 19300 14430 19310 14890
rect 19250 14350 19310 14430
rect 19360 14890 19420 14910
rect 19360 14430 19370 14890
rect 19410 14430 19420 14890
rect 19360 14410 19420 14430
rect 19470 14890 19530 14910
rect 19470 14430 19480 14890
rect 19520 14430 19530 14890
rect 19470 14350 19530 14430
rect 19580 14890 19640 14910
rect 19580 14430 19590 14890
rect 19630 14430 19640 14890
rect 19580 14410 19640 14430
rect 19690 14890 19750 14910
rect 19690 14430 19700 14890
rect 19740 14430 19750 14890
rect 19690 14350 19750 14430
rect 19800 14890 19860 14910
rect 19800 14430 19810 14890
rect 19850 14430 19860 14890
rect 19800 14410 19860 14430
rect 19910 14890 19970 14910
rect 19910 14430 19920 14890
rect 19960 14430 19970 14890
rect 19910 14350 19970 14430
rect 20020 14890 20080 14910
rect 20020 14430 20030 14890
rect 20070 14430 20080 14890
rect 20020 14410 20080 14430
rect 20130 14890 20190 14910
rect 20130 14430 20140 14890
rect 20180 14430 20190 14890
rect 20130 14350 20190 14430
rect 20240 14890 20300 14910
rect 20240 14430 20250 14890
rect 20290 14430 20300 14890
rect 20240 14410 20300 14430
rect 20350 14890 20410 14910
rect 20350 14430 20360 14890
rect 20400 14430 20410 14890
rect 20350 14350 20410 14430
rect 20460 14890 20520 14910
rect 20460 14430 20470 14890
rect 20510 14430 20520 14890
rect 20460 14410 20520 14430
rect 20570 14890 20630 14910
rect 20570 14430 20580 14890
rect 20620 14430 20630 14890
rect 20570 14350 20630 14430
rect 20680 14890 20740 14910
rect 20680 14430 20690 14890
rect 20730 14430 20740 14890
rect 20680 14410 20740 14430
rect 20790 14890 20850 14910
rect 20790 14430 20800 14890
rect 20840 14430 20850 14890
rect 20790 14350 20850 14430
rect 20900 14890 20960 14960
rect 20900 14430 20910 14890
rect 20950 14430 20960 14890
rect 20900 14410 20960 14430
rect 9670 14340 21120 14350
rect 9670 14300 9700 14340
rect 9740 14300 9790 14340
rect 9830 14300 9870 14340
rect 9910 14300 9950 14340
rect 9990 14300 10030 14340
rect 10070 14300 10110 14340
rect 10150 14300 10190 14340
rect 10230 14300 10270 14340
rect 10310 14300 10350 14340
rect 10390 14300 10430 14340
rect 10470 14300 10510 14340
rect 10550 14300 10590 14340
rect 10630 14300 10670 14340
rect 10710 14300 10750 14340
rect 10790 14300 10830 14340
rect 10870 14300 10910 14340
rect 10950 14300 10990 14340
rect 11030 14300 11070 14340
rect 11110 14300 11150 14340
rect 11190 14300 11230 14340
rect 11270 14300 11310 14340
rect 11350 14300 11390 14340
rect 11430 14300 11470 14340
rect 11510 14300 11550 14340
rect 11590 14300 11630 14340
rect 11670 14300 11710 14340
rect 11750 14300 11790 14340
rect 11830 14300 11870 14340
rect 11910 14300 11950 14340
rect 11990 14300 12030 14340
rect 12070 14300 12110 14340
rect 12150 14300 12190 14340
rect 12230 14300 12270 14340
rect 12310 14300 12350 14340
rect 12390 14300 12430 14340
rect 12470 14300 12510 14340
rect 12550 14300 12590 14340
rect 12630 14300 12670 14340
rect 12710 14300 12750 14340
rect 12790 14300 12830 14340
rect 12870 14300 12910 14340
rect 12950 14300 12990 14340
rect 13030 14300 13070 14340
rect 13110 14300 13150 14340
rect 13230 14300 13270 14340
rect 13310 14300 13350 14340
rect 13390 14300 13430 14340
rect 13470 14300 13510 14340
rect 13550 14300 13590 14340
rect 13630 14300 13670 14340
rect 13710 14300 13750 14340
rect 13790 14300 13830 14340
rect 13870 14300 13910 14340
rect 13950 14300 13990 14340
rect 14030 14300 14070 14340
rect 14110 14300 14150 14340
rect 14190 14300 14230 14340
rect 14270 14300 14310 14340
rect 14350 14300 14390 14340
rect 14430 14300 14470 14340
rect 14510 14300 14550 14340
rect 14590 14300 14630 14340
rect 14670 14300 14710 14340
rect 14750 14300 14790 14340
rect 14830 14300 14870 14340
rect 14910 14300 14950 14340
rect 14990 14300 15030 14340
rect 15070 14300 15110 14340
rect 15150 14300 15190 14340
rect 15230 14300 15270 14340
rect 15310 14300 15350 14340
rect 15390 14300 15430 14340
rect 15470 14300 15510 14340
rect 15550 14300 15590 14340
rect 15630 14300 15670 14340
rect 15710 14300 15750 14340
rect 15790 14300 15830 14340
rect 15870 14300 15910 14340
rect 15950 14300 15990 14340
rect 16030 14300 16070 14340
rect 16110 14300 16150 14340
rect 16190 14300 16230 14340
rect 16270 14300 16310 14340
rect 16350 14300 16390 14340
rect 16430 14300 16470 14340
rect 16510 14300 16550 14340
rect 16590 14300 16630 14340
rect 16670 14300 16710 14340
rect 16750 14300 16790 14340
rect 16830 14300 16870 14340
rect 16910 14300 16950 14340
rect 16990 14300 17030 14340
rect 17070 14300 17110 14340
rect 17150 14300 17190 14340
rect 17230 14300 17270 14340
rect 17310 14300 17350 14340
rect 17390 14300 17430 14340
rect 17470 14300 17510 14340
rect 17550 14300 17590 14340
rect 17630 14300 17670 14340
rect 17710 14300 17750 14340
rect 17790 14300 17830 14340
rect 17870 14300 17910 14340
rect 17950 14300 17990 14340
rect 18030 14300 18070 14340
rect 18110 14300 18150 14340
rect 18190 14300 18230 14340
rect 18270 14300 18310 14340
rect 18350 14300 18390 14340
rect 18430 14300 18470 14340
rect 18510 14300 18550 14340
rect 18590 14300 18630 14340
rect 18670 14300 18710 14340
rect 18750 14300 18790 14340
rect 18830 14300 18870 14340
rect 18910 14300 18950 14340
rect 18990 14300 19030 14340
rect 19070 14300 19110 14340
rect 19150 14300 19190 14340
rect 19230 14300 19270 14340
rect 19310 14300 19350 14340
rect 19390 14300 19430 14340
rect 19470 14300 19510 14340
rect 19550 14300 19590 14340
rect 19630 14300 19670 14340
rect 19710 14300 19750 14340
rect 19790 14300 19830 14340
rect 19870 14300 19910 14340
rect 19950 14300 19990 14340
rect 20030 14300 20070 14340
rect 20110 14300 20150 14340
rect 20190 14300 20230 14340
rect 20270 14300 20310 14340
rect 20350 14300 20390 14340
rect 20430 14300 20470 14340
rect 20510 14300 20550 14340
rect 20590 14300 20630 14340
rect 20670 14300 20710 14340
rect 20750 14300 20790 14340
rect 20830 14300 20870 14340
rect 20910 14300 20950 14340
rect 20990 14300 21030 14340
rect 21070 14300 21120 14340
rect 9670 14290 21120 14300
rect 7280 13370 21110 13380
rect 7280 13330 7320 13370
rect 7360 13330 7400 13370
rect 7440 13330 7480 13370
rect 7520 13330 7560 13370
rect 7600 13330 7640 13370
rect 7680 13330 7720 13370
rect 7760 13330 7800 13370
rect 7840 13330 7880 13370
rect 7920 13330 7960 13370
rect 8000 13330 8040 13370
rect 8080 13330 8120 13370
rect 8160 13330 8200 13370
rect 8240 13330 8280 13370
rect 8320 13330 8360 13370
rect 8400 13330 8440 13370
rect 8480 13330 8520 13370
rect 8560 13330 8600 13370
rect 8640 13330 8680 13370
rect 8720 13330 8760 13370
rect 8800 13330 8840 13370
rect 8880 13330 8920 13370
rect 8960 13330 9000 13370
rect 9040 13330 9080 13370
rect 9120 13330 9160 13370
rect 9200 13330 9240 13370
rect 9280 13330 9320 13370
rect 9360 13330 9400 13370
rect 9440 13330 9480 13370
rect 9520 13330 9560 13370
rect 9600 13330 9640 13370
rect 9680 13330 9720 13370
rect 9760 13330 9800 13370
rect 9840 13330 9890 13370
rect 9930 13330 9970 13370
rect 10010 13330 10050 13370
rect 10090 13330 10130 13370
rect 10170 13330 10210 13370
rect 10250 13330 10290 13370
rect 10330 13330 10370 13370
rect 10410 13330 10450 13370
rect 10490 13330 10530 13370
rect 10570 13330 10610 13370
rect 10650 13330 10690 13370
rect 10730 13330 10770 13370
rect 10810 13330 10850 13370
rect 10890 13330 10930 13370
rect 10970 13330 11010 13370
rect 11050 13330 11090 13370
rect 11130 13330 11170 13370
rect 11210 13330 11250 13370
rect 11290 13330 11330 13370
rect 11370 13330 11410 13370
rect 11450 13330 11490 13370
rect 11530 13330 11570 13370
rect 11610 13330 11650 13370
rect 11690 13330 11730 13370
rect 11770 13330 11810 13370
rect 11850 13330 11890 13370
rect 11930 13330 11970 13370
rect 12010 13330 12050 13370
rect 12090 13330 12130 13370
rect 12170 13330 12210 13370
rect 12250 13330 12290 13370
rect 12330 13330 12370 13370
rect 12410 13330 12450 13370
rect 12490 13330 12530 13370
rect 12570 13330 12610 13370
rect 12650 13330 12690 13370
rect 12730 13330 12770 13370
rect 12810 13330 12850 13370
rect 12890 13330 12930 13370
rect 12970 13330 13010 13370
rect 13050 13330 13090 13370
rect 13130 13330 13170 13370
rect 13210 13330 13250 13370
rect 13290 13330 13330 13370
rect 13400 13330 13440 13370
rect 13480 13330 13520 13370
rect 13560 13330 13600 13370
rect 13640 13330 13680 13370
rect 13720 13330 13760 13370
rect 13800 13330 13840 13370
rect 13880 13330 13920 13370
rect 13960 13330 14000 13370
rect 14040 13330 14080 13370
rect 14120 13330 14160 13370
rect 14200 13330 14240 13370
rect 14280 13330 14320 13370
rect 14360 13330 14400 13370
rect 14440 13330 14480 13370
rect 14520 13330 14560 13370
rect 14600 13330 14640 13370
rect 14680 13330 14720 13370
rect 14760 13330 14800 13370
rect 14840 13330 14880 13370
rect 14920 13330 14960 13370
rect 15000 13330 15040 13370
rect 15080 13330 15120 13370
rect 15160 13330 15200 13370
rect 15240 13330 15280 13370
rect 15320 13330 15360 13370
rect 15400 13330 15440 13370
rect 15480 13330 15520 13370
rect 15560 13330 15600 13370
rect 15640 13330 15680 13370
rect 15720 13330 15760 13370
rect 15800 13330 15840 13370
rect 15880 13330 15920 13370
rect 15960 13330 16000 13370
rect 16040 13330 16080 13370
rect 16120 13330 16160 13370
rect 16200 13330 16240 13370
rect 16280 13330 16320 13370
rect 16360 13330 16400 13370
rect 16440 13330 16480 13370
rect 16520 13330 16560 13370
rect 16600 13330 16640 13370
rect 16680 13330 16720 13370
rect 16760 13330 16800 13370
rect 16840 13330 16880 13370
rect 16920 13330 16960 13370
rect 17000 13330 17040 13370
rect 17080 13330 17120 13370
rect 17160 13330 17200 13370
rect 17240 13330 17280 13370
rect 17320 13330 17360 13370
rect 17400 13330 17440 13370
rect 17480 13330 17520 13370
rect 17560 13330 17600 13370
rect 17640 13330 17680 13370
rect 17720 13330 17760 13370
rect 17800 13330 17840 13370
rect 17880 13330 17920 13370
rect 17960 13330 18000 13370
rect 18040 13330 18080 13370
rect 18120 13330 18160 13370
rect 18200 13330 18240 13370
rect 18280 13330 18320 13370
rect 18360 13330 18400 13370
rect 18440 13330 18480 13370
rect 18520 13330 18560 13370
rect 18600 13330 18640 13370
rect 18680 13330 18720 13370
rect 18760 13330 18800 13370
rect 18840 13330 18880 13370
rect 18920 13330 18960 13370
rect 19000 13330 19040 13370
rect 19080 13330 19120 13370
rect 19160 13330 19200 13370
rect 19240 13330 19280 13370
rect 19320 13330 19360 13370
rect 19400 13330 19440 13370
rect 19480 13330 19520 13370
rect 19560 13330 19600 13370
rect 19640 13330 19680 13370
rect 19720 13330 19760 13370
rect 19800 13330 19840 13370
rect 19880 13330 19920 13370
rect 19960 13330 20000 13370
rect 20040 13330 20080 13370
rect 20120 13330 20160 13370
rect 20200 13330 20240 13370
rect 20280 13330 20320 13370
rect 20360 13330 20400 13370
rect 20440 13330 20480 13370
rect 20520 13330 20560 13370
rect 20600 13330 20640 13370
rect 20680 13330 20720 13370
rect 20760 13330 20800 13370
rect 20840 13330 20880 13370
rect 20920 13330 20960 13370
rect 21000 13330 21040 13370
rect 21080 13330 21110 13370
rect 7280 13320 21110 13330
rect 7280 13240 7340 13320
rect 7280 12780 7290 13240
rect 7330 12780 7340 13240
rect 7280 12760 7340 12780
rect 7390 13240 7450 13260
rect 7390 12780 7400 13240
rect 7440 12780 7450 13240
rect 7390 12720 7450 12780
rect 7500 13240 7560 13320
rect 7500 12780 7510 13240
rect 7550 12780 7560 13240
rect 7500 12760 7560 12780
rect 7910 13240 7970 13320
rect 7910 12780 7920 13240
rect 7960 12780 7970 13240
rect 7910 12760 7970 12780
rect 8040 13240 8100 13260
rect 8040 12780 8050 13240
rect 8090 12780 8100 13240
rect 8040 12720 8100 12780
rect 8170 13240 8230 13320
rect 8170 12780 8180 13240
rect 8220 12780 8230 13240
rect 8170 12760 8230 12780
rect 8550 13240 8610 13320
rect 8550 12780 8560 13240
rect 8600 12780 8610 13240
rect 8550 12760 8610 12780
rect 8680 13240 8740 13260
rect 8680 12780 8690 13240
rect 8730 12780 8740 13240
rect 8680 12720 8740 12780
rect 8810 13240 8870 13320
rect 8810 12780 8820 13240
rect 8860 12780 8870 13240
rect 8810 12760 8870 12780
rect 8930 13240 8990 13320
rect 8930 12780 8940 13240
rect 8980 12780 8990 13240
rect 8930 12760 8990 12780
rect 9040 13240 9100 13260
rect 9040 12780 9050 13240
rect 9090 12780 9100 13240
rect 9040 12720 9100 12780
rect 9190 13240 9250 13320
rect 9190 12780 9200 13240
rect 9240 12780 9250 13240
rect 9190 12760 9250 12780
rect 9300 13240 9360 13260
rect 9300 12780 9310 13240
rect 9350 12780 9360 13240
rect 9300 12720 9360 12780
rect 9440 13240 9500 13320
rect 9440 12780 9450 13240
rect 9490 12780 9500 13240
rect 9440 12760 9500 12780
rect 9550 13240 9610 13260
rect 9550 12780 9560 13240
rect 9600 12780 9610 13240
rect 9860 13240 9920 13320
rect 9550 12720 9610 12780
rect 9860 12780 9870 13240
rect 9910 12780 9920 13240
rect 9860 12760 9920 12780
rect 9970 13240 10030 13260
rect 9970 12780 9980 13240
rect 10020 12780 10030 13240
rect 9970 12720 10030 12780
rect 10080 13240 10140 13320
rect 10080 12780 10090 13240
rect 10130 12780 10140 13240
rect 10080 12760 10140 12780
rect 10510 13240 10570 13320
rect 10510 12780 10520 13240
rect 10560 12780 10570 13240
rect 10510 12760 10570 12780
rect 10640 13240 10700 13260
rect 10640 12780 10650 13240
rect 10690 12780 10700 13240
rect 10640 12720 10700 12780
rect 10770 13240 10830 13320
rect 10770 12780 10780 13240
rect 10820 12780 10830 13240
rect 10770 12760 10830 12780
rect 11000 13240 11060 13320
rect 11000 12780 11010 13240
rect 11050 12780 11060 13240
rect 11000 12760 11060 12780
rect 11110 13240 11170 13260
rect 11110 12780 11120 13240
rect 11160 12780 11170 13240
rect 11110 12720 11170 12780
rect 11220 13240 11280 13320
rect 11220 12780 11230 13240
rect 11270 12780 11280 13240
rect 11220 12760 11280 12780
rect 11500 13240 11560 13320
rect 11500 12780 11510 13240
rect 11550 12780 11560 13240
rect 11500 12760 11560 12780
rect 11630 13240 11690 13260
rect 11630 12780 11640 13240
rect 11680 12780 11690 13240
rect 11630 12720 11690 12780
rect 11760 13240 11820 13320
rect 11760 12780 11770 13240
rect 11810 12780 11820 13240
rect 11760 12760 11820 12780
rect 11990 13240 12050 13320
rect 11990 12780 12000 13240
rect 12040 12780 12050 13240
rect 11990 12760 12050 12780
rect 12100 13240 12160 13260
rect 12100 12780 12110 13240
rect 12150 12780 12160 13240
rect 12100 12720 12160 12780
rect 12210 13240 12270 13320
rect 12210 12780 12220 13240
rect 12260 12780 12270 13240
rect 12210 12760 12270 12780
rect 12500 13240 12560 13320
rect 12500 12780 12510 13240
rect 12550 12780 12560 13240
rect 12500 12760 12560 12780
rect 12630 13240 12690 13260
rect 12630 12780 12640 13240
rect 12680 12780 12690 13240
rect 12630 12720 12690 12780
rect 12760 13240 12820 13320
rect 12760 12780 12770 13240
rect 12810 12780 12820 13240
rect 12760 12760 12820 12780
rect 12990 13240 13050 13320
rect 12990 12780 13000 13240
rect 13040 12780 13050 13240
rect 12990 12760 13050 12780
rect 13100 13240 13160 13260
rect 13100 12780 13110 13240
rect 13150 12780 13160 13240
rect 13100 12720 13160 12780
rect 13210 13240 13270 13320
rect 13210 12780 13220 13240
rect 13260 12780 13270 13240
rect 13210 12760 13270 12780
rect 13340 13240 13400 13320
rect 13340 12780 13350 13240
rect 13390 12780 13400 13240
rect 13340 12760 13400 12780
rect 13450 13240 13510 13260
rect 13450 12780 13460 13240
rect 13500 12780 13510 13240
rect 7250 12710 7350 12720
rect 7250 12650 7270 12710
rect 7330 12650 7350 12710
rect 7250 12640 7350 12650
rect 7390 12710 7870 12720
rect 7390 12700 7700 12710
rect 7390 12660 7570 12700
rect 7610 12660 7700 12700
rect 7390 12650 7700 12660
rect 7760 12700 7870 12710
rect 7760 12660 7820 12700
rect 7860 12660 7870 12700
rect 8040 12710 8380 12720
rect 8040 12670 8320 12710
rect 8360 12670 8380 12710
rect 8040 12660 8380 12670
rect 8550 12690 8620 12710
rect 7760 12650 7870 12660
rect 7390 12640 7870 12650
rect 7280 12300 7340 12320
rect 7280 12140 7290 12300
rect 7330 12140 7340 12300
rect 7280 12010 7340 12140
rect 7390 12300 7450 12640
rect 8070 12600 8130 12620
rect 8070 12560 8080 12600
rect 8120 12560 8130 12600
rect 8070 12540 8130 12560
rect 7910 12500 7970 12520
rect 7390 12140 7400 12300
rect 7440 12140 7450 12300
rect 7390 12120 7450 12140
rect 7500 12300 7560 12320
rect 7500 12140 7510 12300
rect 7550 12140 7560 12300
rect 7500 12010 7560 12140
rect 7910 12140 7920 12500
rect 7960 12140 7970 12500
rect 7910 12010 7970 12140
rect 8170 12500 8230 12660
rect 8550 12650 8570 12690
rect 8610 12650 8620 12690
rect 8550 12630 8620 12650
rect 8680 12700 9000 12720
rect 8680 12660 8870 12700
rect 8910 12660 8950 12700
rect 8990 12660 9000 12700
rect 8680 12640 9000 12660
rect 9040 12700 9260 12720
rect 9040 12660 9070 12700
rect 9110 12660 9210 12700
rect 9250 12660 9260 12700
rect 9040 12640 9260 12660
rect 9300 12700 9510 12720
rect 9300 12660 9330 12700
rect 9370 12660 9460 12700
rect 9500 12660 9510 12700
rect 9300 12640 9510 12660
rect 9550 12700 9630 12720
rect 9550 12660 9580 12700
rect 9620 12660 9630 12700
rect 9840 12710 9930 12720
rect 9840 12670 9860 12710
rect 9900 12670 9930 12710
rect 9840 12660 9930 12670
rect 9970 12710 10220 12720
rect 9970 12670 10160 12710
rect 10200 12670 10220 12710
rect 9970 12660 10220 12670
rect 10410 12700 10470 12720
rect 10410 12660 10420 12700
rect 10460 12660 10470 12700
rect 10640 12710 11070 12720
rect 10640 12670 10920 12710
rect 10960 12670 11000 12710
rect 11040 12670 11070 12710
rect 10640 12660 11070 12670
rect 11110 12710 11350 12720
rect 11110 12670 11300 12710
rect 11340 12670 11350 12710
rect 11110 12660 11350 12670
rect 11400 12700 11460 12720
rect 11400 12660 11410 12700
rect 11450 12660 11460 12700
rect 11630 12710 12060 12720
rect 11630 12670 11910 12710
rect 11950 12670 11990 12710
rect 12030 12670 12060 12710
rect 11630 12660 12060 12670
rect 12100 12710 12340 12720
rect 12100 12670 12290 12710
rect 12330 12670 12340 12710
rect 12100 12660 12340 12670
rect 12400 12700 12460 12720
rect 12400 12660 12410 12700
rect 12450 12660 12460 12700
rect 12630 12710 13060 12720
rect 12630 12670 12910 12710
rect 12950 12670 12990 12710
rect 13030 12670 13060 12710
rect 12630 12660 13060 12670
rect 13100 12700 13410 12720
rect 13100 12660 13280 12700
rect 13320 12660 13360 12700
rect 13400 12660 13410 12700
rect 9550 12640 9630 12660
rect 8700 12580 8770 12600
rect 8700 12540 8720 12580
rect 8760 12540 8770 12580
rect 8700 12520 8770 12540
rect 8170 12140 8180 12500
rect 8220 12140 8230 12500
rect 8170 12120 8230 12140
rect 8550 12460 8610 12480
rect 8550 12100 8560 12460
rect 8600 12100 8610 12460
rect 8550 12010 8610 12100
rect 8680 12460 8740 12480
rect 8680 12100 8690 12460
rect 8730 12100 8740 12460
rect 8680 12080 8740 12100
rect 8810 12460 8870 12640
rect 8810 12100 8820 12460
rect 8860 12100 8870 12460
rect 8810 12080 8870 12100
rect 8930 12570 8990 12590
rect 8930 12410 8940 12570
rect 8980 12410 8990 12570
rect 8930 12350 8990 12410
rect 9040 12570 9100 12640
rect 9040 12410 9050 12570
rect 9090 12410 9100 12570
rect 9040 12390 9100 12410
rect 9190 12570 9250 12590
rect 9190 12410 9200 12570
rect 9240 12410 9250 12570
rect 9190 12350 9250 12410
rect 9300 12570 9360 12640
rect 9300 12410 9310 12570
rect 9350 12410 9360 12570
rect 9300 12390 9360 12410
rect 9440 12570 9500 12590
rect 9440 12410 9450 12570
rect 9490 12410 9500 12570
rect 9440 12350 9500 12410
rect 9550 12570 9610 12640
rect 9550 12410 9560 12570
rect 9600 12410 9610 12570
rect 9550 12390 9610 12410
rect 8930 12290 9500 12350
rect 9860 12300 9920 12320
rect 8930 12010 8990 12290
rect 9860 12140 9870 12300
rect 9910 12140 9920 12300
rect 9860 12060 9920 12140
rect 9970 12300 10030 12660
rect 10410 12640 10470 12660
rect 10670 12600 10730 12620
rect 10670 12560 10680 12600
rect 10720 12560 10730 12600
rect 10670 12540 10730 12560
rect 10510 12500 10570 12520
rect 9970 12140 9980 12300
rect 10020 12140 10030 12300
rect 9970 12120 10030 12140
rect 10080 12300 10140 12320
rect 10080 12140 10090 12300
rect 10130 12140 10140 12300
rect 10080 12060 10140 12140
rect 10510 12140 10520 12500
rect 10560 12140 10570 12500
rect 10510 12060 10570 12140
rect 10770 12500 10830 12660
rect 10770 12140 10780 12500
rect 10820 12140 10830 12500
rect 10770 12120 10830 12140
rect 11000 12300 11060 12320
rect 11000 12140 11010 12300
rect 11050 12140 11060 12300
rect 11000 12060 11060 12140
rect 11110 12300 11170 12660
rect 11400 12640 11460 12660
rect 11660 12600 11720 12620
rect 11660 12560 11670 12600
rect 11710 12560 11720 12600
rect 11660 12540 11720 12560
rect 11500 12500 11560 12520
rect 11110 12140 11120 12300
rect 11160 12140 11170 12300
rect 11110 12120 11170 12140
rect 11220 12300 11280 12320
rect 11220 12140 11230 12300
rect 11270 12140 11280 12300
rect 11220 12060 11280 12140
rect 11500 12140 11510 12500
rect 11550 12140 11560 12500
rect 11500 12060 11560 12140
rect 11760 12500 11820 12660
rect 11760 12140 11770 12500
rect 11810 12140 11820 12500
rect 11760 12120 11820 12140
rect 11990 12300 12050 12320
rect 11990 12140 12000 12300
rect 12040 12140 12050 12300
rect 11990 12060 12050 12140
rect 12100 12300 12160 12660
rect 12400 12640 12460 12660
rect 12660 12600 12720 12620
rect 12660 12560 12670 12600
rect 12710 12560 12720 12600
rect 12660 12540 12720 12560
rect 12500 12500 12560 12520
rect 12100 12140 12110 12300
rect 12150 12140 12160 12300
rect 12100 12120 12160 12140
rect 12210 12300 12270 12320
rect 12210 12140 12220 12300
rect 12260 12140 12270 12300
rect 12210 12060 12270 12140
rect 12500 12140 12510 12500
rect 12550 12140 12560 12500
rect 12500 12060 12560 12140
rect 12760 12500 12820 12660
rect 12760 12140 12770 12500
rect 12810 12140 12820 12500
rect 13100 12640 13410 12660
rect 13450 12700 13510 12780
rect 13570 13240 13630 13260
rect 13570 12780 13580 13240
rect 13620 12780 13630 13240
rect 13570 12760 13630 12780
rect 13680 13240 13740 13320
rect 13680 12780 13690 13240
rect 13730 12780 13740 13240
rect 13680 12760 13740 12780
rect 13790 13240 13850 13260
rect 13790 12780 13800 13240
rect 13840 12780 13850 13240
rect 13450 12660 13460 12700
rect 13500 12660 13510 12700
rect 12760 12120 12820 12140
rect 12990 12300 13050 12320
rect 12990 12140 13000 12300
rect 13040 12140 13050 12300
rect 12990 12060 13050 12140
rect 13100 12300 13160 12640
rect 13340 12580 13400 12600
rect 13340 12420 13350 12580
rect 13390 12420 13400 12580
rect 13100 12140 13110 12300
rect 13150 12140 13160 12300
rect 13100 12120 13160 12140
rect 13210 12300 13270 12320
rect 13210 12140 13220 12300
rect 13260 12140 13270 12300
rect 13210 12060 13270 12140
rect 13340 12060 13400 12420
rect 13450 12580 13510 12660
rect 13580 12700 13640 12720
rect 13580 12660 13590 12700
rect 13630 12660 13640 12700
rect 13580 12640 13640 12660
rect 13790 12700 13850 12780
rect 13910 13240 13970 13260
rect 13910 12780 13920 13240
rect 13960 12780 13970 13240
rect 13910 12760 13970 12780
rect 14020 13240 14080 13320
rect 14020 12780 14030 13240
rect 14070 12780 14080 13240
rect 14020 12760 14080 12780
rect 14130 13240 14190 13260
rect 14130 12780 14140 13240
rect 14180 12780 14190 13240
rect 14130 12760 14190 12780
rect 14240 13240 14300 13320
rect 14240 12780 14250 13240
rect 14290 12780 14300 13240
rect 14240 12760 14300 12780
rect 14350 13240 14410 13260
rect 14350 12780 14360 13240
rect 14400 12780 14410 13240
rect 13790 12660 13800 12700
rect 13840 12660 13850 12700
rect 13450 12420 13460 12580
rect 13500 12420 13510 12580
rect 13450 12400 13510 12420
rect 13570 12580 13630 12600
rect 13570 12420 13580 12580
rect 13620 12420 13630 12580
rect 13570 12400 13630 12420
rect 13680 12580 13740 12600
rect 13680 12420 13690 12580
rect 13730 12420 13740 12580
rect 13680 12060 13740 12420
rect 13790 12580 13850 12660
rect 13920 12700 13980 12720
rect 13920 12660 13930 12700
rect 13970 12660 13980 12700
rect 13920 12640 13980 12660
rect 14350 12700 14410 12780
rect 14470 13240 14530 13260
rect 14470 12780 14480 13240
rect 14520 12780 14530 13240
rect 14470 12760 14530 12780
rect 14580 13240 14640 13320
rect 14580 12780 14590 13240
rect 14630 12780 14640 13240
rect 14580 12760 14640 12780
rect 14690 13240 14750 13260
rect 14690 12780 14700 13240
rect 14740 12780 14750 13240
rect 14690 12760 14750 12780
rect 14800 13240 14860 13320
rect 14800 12780 14810 13240
rect 14850 12780 14860 13240
rect 14800 12760 14860 12780
rect 14910 13240 14970 13260
rect 14910 12780 14920 13240
rect 14960 12780 14970 13240
rect 14910 12760 14970 12780
rect 15020 13240 15080 13320
rect 15020 12780 15030 13240
rect 15070 12780 15080 13240
rect 15020 12760 15080 12780
rect 15130 13240 15190 13260
rect 15130 12780 15140 13240
rect 15180 12780 15190 13240
rect 15130 12760 15190 12780
rect 15240 13240 15300 13320
rect 15240 12780 15250 13240
rect 15290 12780 15300 13240
rect 15240 12760 15300 12780
rect 15350 13240 15410 13260
rect 15350 12780 15360 13240
rect 15400 12780 15410 13240
rect 14350 12660 14360 12700
rect 14400 12660 14410 12700
rect 13790 12420 13800 12580
rect 13840 12420 13850 12580
rect 13790 12400 13850 12420
rect 13910 12580 13970 12600
rect 13910 12420 13920 12580
rect 13960 12420 13970 12580
rect 13910 12400 13970 12420
rect 14020 12580 14080 12600
rect 14020 12420 14030 12580
rect 14070 12420 14080 12580
rect 14020 12060 14080 12420
rect 14130 12580 14190 12600
rect 14130 12420 14140 12580
rect 14180 12420 14190 12580
rect 14130 12400 14190 12420
rect 14240 12580 14300 12600
rect 14240 12420 14250 12580
rect 14290 12420 14300 12580
rect 14240 12060 14300 12420
rect 14350 12580 14410 12660
rect 14480 12700 14540 12720
rect 14480 12660 14490 12700
rect 14530 12660 14540 12700
rect 14480 12640 14540 12660
rect 15350 12700 15410 12780
rect 15530 13240 15590 13260
rect 15530 12780 15540 13240
rect 15580 12780 15590 13240
rect 15530 12760 15590 12780
rect 15640 13240 15700 13320
rect 15640 12780 15650 13240
rect 15690 12780 15700 13240
rect 15640 12760 15700 12780
rect 15750 13240 15810 13260
rect 15750 12780 15760 13240
rect 15800 12780 15810 13240
rect 15750 12760 15810 12780
rect 15860 13240 15920 13320
rect 15860 12780 15870 13240
rect 15910 12780 15920 13240
rect 15860 12760 15920 12780
rect 15970 13240 16030 13260
rect 15970 12780 15980 13240
rect 16020 12780 16030 13240
rect 15970 12760 16030 12780
rect 16080 13240 16140 13320
rect 16080 12780 16090 13240
rect 16130 12780 16140 13240
rect 16080 12760 16140 12780
rect 16190 13240 16250 13260
rect 16190 12780 16200 13240
rect 16240 12780 16250 13240
rect 16190 12760 16250 12780
rect 16300 13240 16360 13320
rect 16300 12780 16310 13240
rect 16350 12780 16360 13240
rect 16300 12760 16360 12780
rect 16410 13240 16470 13260
rect 16410 12780 16420 13240
rect 16460 12780 16470 13240
rect 16410 12760 16470 12780
rect 16520 13240 16580 13320
rect 16520 12780 16530 13240
rect 16570 12780 16580 13240
rect 16520 12760 16580 12780
rect 16630 13240 16690 13260
rect 16630 12780 16640 13240
rect 16680 12780 16690 13240
rect 16630 12760 16690 12780
rect 16740 13240 16800 13320
rect 16740 12780 16750 13240
rect 16790 12780 16800 13240
rect 16740 12760 16800 12780
rect 16850 13240 16910 13260
rect 16850 12780 16860 13240
rect 16900 12780 16910 13240
rect 16850 12760 16910 12780
rect 16960 13240 17020 13320
rect 16960 12780 16970 13240
rect 17010 12780 17020 13240
rect 16960 12760 17020 12780
rect 17070 13240 17130 13260
rect 17070 12780 17080 13240
rect 17120 12780 17130 13240
rect 17070 12760 17130 12780
rect 17180 13240 17240 13320
rect 17180 12780 17190 13240
rect 17230 12780 17240 13240
rect 17180 12760 17240 12780
rect 17290 13240 17350 13260
rect 17290 12780 17300 13240
rect 17340 12780 17350 13240
rect 15350 12660 15360 12700
rect 15400 12660 15410 12700
rect 14350 12420 14360 12580
rect 14400 12420 14410 12580
rect 14350 12400 14410 12420
rect 14470 12580 14530 12600
rect 14470 12420 14480 12580
rect 14520 12420 14530 12580
rect 14470 12400 14530 12420
rect 14580 12580 14640 12600
rect 14580 12420 14590 12580
rect 14630 12420 14640 12580
rect 14580 12060 14640 12420
rect 14690 12580 14750 12600
rect 14690 12420 14700 12580
rect 14740 12420 14750 12580
rect 14690 12400 14750 12420
rect 14800 12580 14860 12600
rect 14800 12420 14810 12580
rect 14850 12420 14860 12580
rect 14800 12060 14860 12420
rect 14910 12580 14970 12600
rect 14910 12420 14920 12580
rect 14960 12420 14970 12580
rect 14910 12400 14970 12420
rect 15020 12580 15080 12600
rect 15020 12420 15030 12580
rect 15070 12420 15080 12580
rect 15020 12060 15080 12420
rect 15130 12580 15190 12600
rect 15130 12420 15140 12580
rect 15180 12420 15190 12580
rect 15130 12400 15190 12420
rect 15240 12580 15300 12600
rect 15240 12420 15250 12580
rect 15290 12420 15300 12580
rect 15240 12060 15300 12420
rect 15350 12580 15410 12660
rect 15540 12700 15600 12720
rect 15540 12660 15550 12700
rect 15590 12660 15600 12700
rect 15540 12640 15600 12660
rect 17290 12710 17350 12780
rect 17480 13240 17540 13260
rect 17480 12780 17490 13240
rect 17530 12780 17540 13240
rect 17480 12760 17540 12780
rect 17590 13240 17650 13320
rect 17590 12780 17600 13240
rect 17640 12780 17650 13240
rect 17590 12760 17650 12780
rect 17700 13240 17760 13260
rect 17700 12780 17710 13240
rect 17750 12780 17760 13240
rect 17700 12760 17760 12780
rect 17810 13240 17870 13320
rect 17810 12780 17820 13240
rect 17860 12780 17870 13240
rect 17810 12760 17870 12780
rect 17920 13240 17980 13260
rect 17920 12780 17930 13240
rect 17970 12780 17980 13240
rect 17920 12760 17980 12780
rect 18030 13240 18090 13320
rect 18030 12780 18040 13240
rect 18080 12780 18090 13240
rect 18030 12760 18090 12780
rect 18140 13240 18200 13260
rect 18140 12780 18150 13240
rect 18190 12780 18200 13240
rect 18140 12760 18200 12780
rect 18250 13240 18310 13320
rect 18250 12780 18260 13240
rect 18300 12780 18310 13240
rect 18250 12760 18310 12780
rect 18360 13240 18420 13260
rect 18360 12780 18370 13240
rect 18410 12780 18420 13240
rect 18360 12760 18420 12780
rect 18470 13240 18530 13320
rect 18470 12780 18480 13240
rect 18520 12780 18530 13240
rect 18470 12760 18530 12780
rect 18580 13240 18640 13260
rect 18580 12780 18590 13240
rect 18630 12780 18640 13240
rect 18580 12760 18640 12780
rect 18690 13240 18750 13320
rect 18690 12780 18700 13240
rect 18740 12780 18750 13240
rect 18690 12760 18750 12780
rect 18800 13240 18860 13260
rect 18800 12780 18810 13240
rect 18850 12780 18860 13240
rect 18800 12760 18860 12780
rect 18910 13240 18970 13320
rect 18910 12780 18920 13240
rect 18960 12780 18970 13240
rect 18910 12760 18970 12780
rect 19020 13240 19080 13260
rect 19020 12780 19030 13240
rect 19070 12780 19080 13240
rect 19020 12760 19080 12780
rect 19130 13240 19190 13320
rect 19130 12780 19140 13240
rect 19180 12780 19190 13240
rect 19130 12760 19190 12780
rect 19240 13240 19300 13260
rect 19240 12780 19250 13240
rect 19290 12780 19300 13240
rect 19240 12760 19300 12780
rect 19350 13240 19410 13320
rect 19350 12780 19360 13240
rect 19400 12780 19410 13240
rect 19350 12760 19410 12780
rect 19460 13240 19520 13260
rect 19460 12780 19470 13240
rect 19510 12780 19520 13240
rect 19460 12760 19520 12780
rect 19570 13240 19630 13320
rect 19570 12780 19580 13240
rect 19620 12780 19630 13240
rect 19570 12760 19630 12780
rect 19680 13240 19740 13260
rect 19680 12780 19690 13240
rect 19730 12780 19740 13240
rect 19680 12760 19740 12780
rect 19790 13240 19850 13320
rect 19790 12780 19800 13240
rect 19840 12780 19850 13240
rect 19790 12760 19850 12780
rect 19900 13240 19960 13260
rect 19900 12780 19910 13240
rect 19950 12780 19960 13240
rect 19900 12760 19960 12780
rect 20010 13240 20070 13320
rect 20010 12780 20020 13240
rect 20060 12780 20070 13240
rect 20010 12760 20070 12780
rect 20120 13240 20180 13260
rect 20120 12780 20130 13240
rect 20170 12780 20180 13240
rect 20120 12760 20180 12780
rect 20230 13240 20290 13320
rect 20230 12780 20240 13240
rect 20280 12780 20290 13240
rect 20230 12760 20290 12780
rect 20340 13240 20400 13260
rect 20340 12780 20350 13240
rect 20390 12780 20400 13240
rect 20340 12760 20400 12780
rect 20450 13240 20510 13320
rect 20450 12780 20460 13240
rect 20500 12780 20510 13240
rect 20450 12760 20510 12780
rect 20560 13240 20620 13260
rect 20560 12780 20570 13240
rect 20610 12780 20620 13240
rect 20560 12760 20620 12780
rect 20670 13240 20730 13320
rect 20670 12780 20680 13240
rect 20720 12780 20730 13240
rect 20670 12760 20730 12780
rect 20780 13240 20840 13260
rect 20780 12780 20790 13240
rect 20830 12780 20840 13240
rect 20780 12760 20840 12780
rect 20890 13240 20950 13320
rect 20890 12780 20900 13240
rect 20940 12780 20950 13240
rect 20890 12760 20950 12780
rect 21000 13240 21060 13260
rect 21000 12780 21010 13240
rect 21050 12780 21060 13240
rect 17290 12700 17420 12710
rect 17290 12650 17350 12700
rect 17400 12650 17420 12700
rect 17290 12640 17420 12650
rect 17480 12700 17550 12720
rect 17480 12660 17500 12700
rect 17540 12660 17550 12700
rect 17480 12640 17550 12660
rect 21000 12710 21060 12780
rect 21000 12700 21130 12710
rect 21000 12650 21060 12700
rect 21110 12650 21130 12700
rect 21000 12640 21130 12650
rect 15350 12420 15360 12580
rect 15400 12420 15410 12580
rect 15350 12400 15410 12420
rect 15530 12580 15590 12600
rect 15530 12420 15540 12580
rect 15580 12420 15590 12580
rect 15530 12400 15590 12420
rect 15640 12580 15700 12600
rect 15640 12420 15650 12580
rect 15690 12420 15700 12580
rect 15640 12060 15700 12420
rect 15750 12580 15810 12600
rect 15750 12420 15760 12580
rect 15800 12420 15810 12580
rect 15750 12400 15810 12420
rect 15860 12580 15920 12600
rect 15860 12420 15870 12580
rect 15910 12420 15920 12580
rect 15860 12060 15920 12420
rect 15970 12580 16030 12600
rect 15970 12420 15980 12580
rect 16020 12420 16030 12580
rect 15970 12400 16030 12420
rect 16080 12580 16140 12600
rect 16080 12420 16090 12580
rect 16130 12420 16140 12580
rect 16080 12060 16140 12420
rect 16190 12580 16250 12600
rect 16190 12420 16200 12580
rect 16240 12420 16250 12580
rect 16190 12400 16250 12420
rect 16300 12580 16360 12600
rect 16300 12420 16310 12580
rect 16350 12420 16360 12580
rect 16300 12060 16360 12420
rect 16410 12580 16470 12600
rect 16410 12420 16420 12580
rect 16460 12420 16470 12580
rect 16410 12400 16470 12420
rect 16520 12580 16580 12600
rect 16520 12420 16530 12580
rect 16570 12420 16580 12580
rect 16520 12060 16580 12420
rect 16630 12580 16690 12600
rect 16630 12420 16640 12580
rect 16680 12420 16690 12580
rect 16630 12400 16690 12420
rect 16740 12580 16800 12600
rect 16740 12420 16750 12580
rect 16790 12420 16800 12580
rect 16740 12060 16800 12420
rect 16850 12580 16910 12600
rect 16850 12420 16860 12580
rect 16900 12420 16910 12580
rect 16850 12400 16910 12420
rect 16960 12580 17020 12600
rect 16960 12420 16970 12580
rect 17010 12420 17020 12580
rect 16960 12060 17020 12420
rect 17070 12580 17130 12600
rect 17070 12420 17080 12580
rect 17120 12420 17130 12580
rect 17070 12400 17130 12420
rect 17180 12580 17240 12600
rect 17180 12420 17190 12580
rect 17230 12420 17240 12580
rect 17180 12060 17240 12420
rect 17290 12580 17350 12640
rect 17290 12420 17300 12580
rect 17340 12420 17350 12580
rect 17290 12400 17350 12420
rect 17480 12580 17540 12600
rect 17480 12420 17490 12580
rect 17530 12420 17540 12580
rect 17480 12400 17540 12420
rect 17590 12580 17650 12600
rect 17590 12420 17600 12580
rect 17640 12420 17650 12580
rect 17590 12060 17650 12420
rect 17700 12580 17760 12600
rect 17700 12420 17710 12580
rect 17750 12420 17760 12580
rect 17700 12400 17760 12420
rect 17810 12580 17870 12600
rect 17810 12420 17820 12580
rect 17860 12420 17870 12580
rect 17810 12060 17870 12420
rect 17920 12580 17980 12600
rect 17920 12420 17930 12580
rect 17970 12420 17980 12580
rect 17920 12400 17980 12420
rect 18030 12580 18090 12600
rect 18030 12420 18040 12580
rect 18080 12420 18090 12580
rect 18030 12060 18090 12420
rect 18140 12580 18200 12600
rect 18140 12420 18150 12580
rect 18190 12420 18200 12580
rect 18140 12400 18200 12420
rect 18250 12580 18310 12600
rect 18250 12420 18260 12580
rect 18300 12420 18310 12580
rect 18250 12060 18310 12420
rect 18360 12580 18420 12600
rect 18360 12420 18370 12580
rect 18410 12420 18420 12580
rect 18360 12400 18420 12420
rect 18470 12580 18530 12600
rect 18470 12420 18480 12580
rect 18520 12420 18530 12580
rect 18470 12060 18530 12420
rect 18580 12580 18640 12600
rect 18580 12420 18590 12580
rect 18630 12420 18640 12580
rect 18580 12400 18640 12420
rect 18690 12580 18750 12600
rect 18690 12420 18700 12580
rect 18740 12420 18750 12580
rect 18690 12060 18750 12420
rect 18800 12580 18860 12600
rect 18800 12420 18810 12580
rect 18850 12420 18860 12580
rect 18800 12400 18860 12420
rect 18910 12580 18970 12600
rect 18910 12420 18920 12580
rect 18960 12420 18970 12580
rect 18910 12060 18970 12420
rect 19020 12580 19080 12600
rect 19020 12420 19030 12580
rect 19070 12420 19080 12580
rect 19020 12400 19080 12420
rect 19130 12580 19190 12600
rect 19130 12420 19140 12580
rect 19180 12420 19190 12580
rect 19130 12060 19190 12420
rect 19240 12580 19300 12600
rect 19240 12420 19250 12580
rect 19290 12420 19300 12580
rect 19240 12400 19300 12420
rect 19350 12580 19410 12600
rect 19350 12420 19360 12580
rect 19400 12420 19410 12580
rect 19350 12060 19410 12420
rect 19460 12580 19520 12600
rect 19460 12420 19470 12580
rect 19510 12420 19520 12580
rect 19460 12400 19520 12420
rect 19570 12580 19630 12600
rect 19570 12420 19580 12580
rect 19620 12420 19630 12580
rect 19570 12060 19630 12420
rect 19680 12580 19740 12600
rect 19680 12420 19690 12580
rect 19730 12420 19740 12580
rect 19680 12400 19740 12420
rect 19790 12580 19850 12600
rect 19790 12420 19800 12580
rect 19840 12420 19850 12580
rect 19790 12060 19850 12420
rect 19900 12580 19960 12600
rect 19900 12420 19910 12580
rect 19950 12420 19960 12580
rect 19900 12400 19960 12420
rect 20010 12580 20070 12600
rect 20010 12420 20020 12580
rect 20060 12420 20070 12580
rect 20010 12060 20070 12420
rect 20120 12580 20180 12600
rect 20120 12420 20130 12580
rect 20170 12420 20180 12580
rect 20120 12400 20180 12420
rect 20230 12580 20290 12600
rect 20230 12420 20240 12580
rect 20280 12420 20290 12580
rect 20230 12060 20290 12420
rect 20340 12580 20400 12600
rect 20340 12420 20350 12580
rect 20390 12420 20400 12580
rect 20340 12400 20400 12420
rect 20450 12580 20510 12600
rect 20450 12420 20460 12580
rect 20500 12420 20510 12580
rect 20450 12060 20510 12420
rect 20560 12580 20620 12600
rect 20560 12420 20570 12580
rect 20610 12420 20620 12580
rect 20560 12400 20620 12420
rect 20670 12580 20730 12600
rect 20670 12420 20680 12580
rect 20720 12420 20730 12580
rect 20670 12060 20730 12420
rect 20780 12580 20840 12600
rect 20780 12420 20790 12580
rect 20830 12420 20840 12580
rect 20780 12400 20840 12420
rect 20890 12580 20950 12600
rect 20890 12420 20900 12580
rect 20940 12420 20950 12580
rect 20890 12060 20950 12420
rect 21000 12580 21060 12640
rect 21000 12420 21010 12580
rect 21050 12420 21060 12580
rect 21000 12400 21060 12420
rect 9730 12050 21160 12060
rect 9730 12010 9810 12050
rect 9850 12010 9890 12050
rect 9930 12010 9970 12050
rect 10010 12010 10050 12050
rect 10090 12010 10130 12050
rect 10170 12010 10210 12050
rect 10250 12010 10290 12050
rect 10330 12010 10370 12050
rect 10410 12010 10450 12050
rect 10490 12010 10530 12050
rect 10570 12010 10610 12050
rect 10650 12010 10690 12050
rect 10730 12010 10770 12050
rect 10810 12010 10850 12050
rect 10890 12010 10930 12050
rect 10970 12010 11010 12050
rect 11050 12010 11090 12050
rect 11130 12010 11170 12050
rect 11210 12010 11250 12050
rect 11290 12010 11330 12050
rect 11370 12010 11410 12050
rect 11450 12010 11490 12050
rect 11530 12010 11570 12050
rect 11610 12010 11650 12050
rect 11690 12010 11730 12050
rect 11770 12010 11810 12050
rect 11850 12010 11890 12050
rect 11930 12010 11970 12050
rect 12010 12010 12050 12050
rect 12090 12010 12130 12050
rect 12170 12010 12210 12050
rect 12250 12010 12290 12050
rect 12330 12010 12370 12050
rect 12410 12010 12450 12050
rect 12490 12010 12530 12050
rect 12570 12010 12610 12050
rect 12650 12010 12690 12050
rect 12730 12010 12770 12050
rect 12810 12010 12850 12050
rect 12890 12010 12930 12050
rect 12970 12010 13010 12050
rect 13050 12010 13090 12050
rect 13130 12010 13170 12050
rect 13210 12010 13250 12050
rect 13290 12010 13330 12050
rect 13440 12010 13480 12050
rect 13520 12010 13560 12050
rect 13600 12010 13640 12050
rect 13680 12010 13720 12050
rect 13760 12010 13800 12050
rect 13840 12010 13880 12050
rect 13920 12010 13960 12050
rect 14000 12010 14040 12050
rect 14080 12010 14120 12050
rect 14160 12010 14200 12050
rect 14240 12010 14280 12050
rect 14320 12010 14360 12050
rect 14400 12010 14440 12050
rect 14480 12010 14520 12050
rect 14560 12010 14600 12050
rect 14640 12010 14680 12050
rect 14720 12010 14760 12050
rect 14800 12010 14840 12050
rect 14880 12010 14920 12050
rect 14960 12010 15000 12050
rect 15040 12010 15080 12050
rect 15120 12010 15160 12050
rect 15200 12010 15240 12050
rect 15280 12010 15320 12050
rect 15360 12010 15400 12050
rect 15440 12010 15480 12050
rect 15520 12010 15560 12050
rect 15600 12010 15640 12050
rect 15680 12010 15720 12050
rect 15760 12010 15800 12050
rect 15840 12010 15880 12050
rect 15920 12010 15960 12050
rect 16000 12010 16040 12050
rect 16080 12010 16120 12050
rect 16160 12010 16200 12050
rect 16240 12010 16280 12050
rect 16320 12010 16360 12050
rect 16400 12010 16440 12050
rect 16480 12010 16520 12050
rect 16560 12010 16600 12050
rect 16640 12010 16680 12050
rect 16720 12010 16760 12050
rect 16800 12010 16840 12050
rect 16880 12010 16920 12050
rect 16960 12010 17000 12050
rect 17040 12010 17080 12050
rect 17120 12010 17160 12050
rect 17200 12010 17240 12050
rect 17280 12010 17320 12050
rect 17360 12010 17400 12050
rect 17440 12010 17480 12050
rect 17520 12010 17560 12050
rect 17600 12010 17640 12050
rect 17680 12010 17720 12050
rect 17760 12010 17800 12050
rect 17840 12010 17880 12050
rect 17920 12010 17960 12050
rect 18000 12010 18040 12050
rect 18080 12010 18120 12050
rect 18160 12010 18200 12050
rect 18240 12010 18280 12050
rect 18320 12010 18360 12050
rect 18400 12010 18440 12050
rect 18480 12010 18520 12050
rect 18560 12010 18600 12050
rect 18640 12010 18680 12050
rect 18720 12010 18760 12050
rect 18800 12010 18840 12050
rect 18880 12010 18920 12050
rect 18960 12010 19000 12050
rect 19040 12010 19080 12050
rect 19120 12010 19160 12050
rect 19200 12010 19240 12050
rect 19280 12010 19320 12050
rect 19360 12010 19400 12050
rect 19440 12010 19480 12050
rect 19520 12010 19560 12050
rect 19600 12010 19640 12050
rect 19680 12010 19720 12050
rect 19760 12010 19800 12050
rect 19840 12010 19890 12050
rect 19930 12010 19970 12050
rect 20010 12010 20050 12050
rect 20090 12010 20130 12050
rect 20170 12010 20210 12050
rect 20250 12010 20290 12050
rect 20330 12010 20370 12050
rect 20410 12010 20460 12050
rect 20500 12010 20540 12050
rect 20580 12010 20620 12050
rect 20660 12010 20700 12050
rect 20740 12010 20780 12050
rect 20820 12010 20860 12050
rect 20900 12010 20940 12050
rect 20980 12010 21020 12050
rect 21060 12010 21160 12050
rect 7280 12000 21160 12010
rect 7280 11960 7330 12000
rect 7370 11960 7410 12000
rect 7450 11960 7490 12000
rect 7530 11960 7570 12000
rect 7610 11960 7650 12000
rect 7690 11960 7730 12000
rect 7770 11960 7810 12000
rect 7850 11960 7890 12000
rect 7930 11960 7970 12000
rect 8010 11960 8050 12000
rect 8090 11960 8130 12000
rect 8170 11960 8210 12000
rect 8250 11960 8290 12000
rect 8330 11960 8370 12000
rect 8410 11960 8450 12000
rect 8490 11960 8530 12000
rect 8570 11960 8610 12000
rect 8650 11960 8690 12000
rect 8730 11960 8770 12000
rect 8810 11960 8850 12000
rect 8890 11960 8930 12000
rect 8970 11960 9010 12000
rect 9050 11960 9090 12000
rect 9130 11960 9170 12000
rect 9210 11960 9250 12000
rect 9290 11960 9330 12000
rect 9370 11960 9410 12000
rect 9450 11960 9490 12000
rect 9530 11960 9570 12000
rect 9610 11960 9650 12000
rect 9690 11960 9730 12000
rect 9770 11960 9800 12000
rect 7280 11950 9800 11960
rect 7660 11410 8600 11420
rect 7660 11370 7720 11410
rect 7760 11370 7800 11410
rect 7840 11370 7880 11410
rect 7920 11370 7960 11410
rect 8000 11370 8040 11410
rect 8080 11370 8120 11410
rect 8160 11370 8200 11410
rect 8240 11370 8280 11410
rect 8320 11370 8360 11410
rect 8400 11370 8440 11410
rect 8480 11370 8520 11410
rect 8560 11370 8600 11410
rect 7660 11360 8600 11370
rect 7660 11330 7720 11360
rect 7660 11290 7670 11330
rect 7710 11290 7720 11330
rect 7660 11250 7720 11290
rect 7660 11210 7670 11250
rect 7710 11210 7720 11250
rect 7660 11170 7720 11210
rect 7660 11130 7670 11170
rect 7710 11130 7720 11170
rect 7660 11100 7720 11130
rect 7280 11090 7720 11100
rect 7280 11050 7330 11090
rect 7370 11050 7410 11090
rect 7450 11050 7490 11090
rect 7530 11050 7570 11090
rect 7610 11050 7650 11090
rect 7690 11050 7720 11090
rect 7280 11040 7720 11050
rect 7850 11280 7910 11300
rect 7850 11120 7860 11280
rect 7900 11120 7910 11280
rect 7850 11060 7910 11120
rect 7960 11280 8020 11360
rect 7960 11120 7970 11280
rect 8010 11120 8020 11280
rect 7960 11100 8020 11120
rect 8090 11280 8150 11300
rect 8090 11120 8100 11280
rect 8140 11120 8150 11280
rect 8090 11060 8150 11120
rect 8220 11280 8280 11360
rect 8540 11330 8600 11360
rect 8220 11120 8230 11280
rect 8270 11120 8280 11280
rect 8220 11100 8280 11120
rect 8330 11280 8390 11300
rect 8330 11120 8340 11280
rect 8380 11120 8390 11280
rect 8330 11060 8390 11120
rect 7280 10910 7340 11040
rect 7280 10750 7290 10910
rect 7330 10750 7340 10910
rect 7280 10730 7340 10750
rect 7390 10910 7450 10930
rect 7390 10750 7400 10910
rect 7440 10750 7450 10910
rect 7250 10410 7350 10420
rect 7250 10350 7270 10410
rect 7330 10350 7350 10410
rect 7250 10340 7350 10350
rect 7390 10390 7450 10750
rect 7500 10910 7560 11040
rect 7850 11000 8390 11060
rect 8540 11290 8550 11330
rect 8590 11290 8600 11330
rect 8540 11250 8600 11290
rect 8540 11210 8550 11250
rect 8590 11210 8600 11250
rect 8540 11170 8600 11210
rect 8540 11130 8550 11170
rect 8590 11130 8600 11170
rect 8540 11100 8600 11130
rect 8540 11090 9800 11100
rect 8540 11050 8610 11090
rect 8650 11050 8690 11090
rect 8730 11050 8770 11090
rect 8810 11050 8850 11090
rect 8890 11050 8930 11090
rect 8970 11050 9010 11090
rect 9050 11050 9090 11090
rect 9130 11050 9170 11090
rect 9210 11050 9250 11090
rect 9290 11050 9330 11090
rect 9370 11050 9410 11090
rect 9450 11050 9490 11090
rect 9530 11050 9570 11090
rect 9610 11050 9650 11090
rect 9690 11050 9730 11090
rect 9770 11050 9800 11090
rect 8540 11040 21160 11050
rect 7500 10750 7510 10910
rect 7550 10750 7560 10910
rect 8120 10940 8180 10960
rect 8120 10900 8130 10940
rect 8170 10900 8180 10940
rect 8120 10880 8180 10900
rect 8330 10950 8390 11000
rect 8640 10960 8700 11040
rect 8330 10940 8430 10950
rect 8330 10900 8350 10940
rect 8390 10900 8430 10940
rect 8330 10890 8430 10900
rect 7840 10850 7920 10870
rect 7840 10790 7850 10850
rect 7910 10790 7920 10850
rect 7840 10770 7920 10790
rect 8330 10780 8390 10890
rect 7500 10730 7560 10750
rect 8220 10720 8390 10780
rect 7960 10700 8020 10720
rect 7390 10380 7670 10390
rect 7390 10340 7610 10380
rect 7650 10340 7670 10380
rect 7390 10330 7670 10340
rect 7280 10270 7340 10290
rect 7280 9810 7290 10270
rect 7330 9810 7340 10270
rect 7280 9730 7340 9810
rect 7390 10270 7450 10330
rect 7390 9810 7400 10270
rect 7440 9810 7450 10270
rect 7390 9790 7450 9810
rect 7500 10270 7560 10290
rect 7500 9810 7510 10270
rect 7550 9810 7560 10270
rect 7500 9730 7560 9810
rect 7960 9740 7970 10700
rect 8010 9740 8020 10700
rect 7280 9720 7790 9730
rect 7280 9680 7320 9720
rect 7360 9680 7400 9720
rect 7440 9680 7480 9720
rect 7520 9680 7560 9720
rect 7600 9680 7640 9720
rect 7680 9680 7720 9720
rect 7760 9680 7790 9720
rect 7280 9670 7790 9680
rect 7710 9650 7790 9670
rect 7960 9650 8020 9740
rect 8220 10700 8280 10720
rect 8220 9740 8230 10700
rect 8270 9740 8280 10700
rect 8640 10600 8650 10960
rect 8690 10600 8700 10960
rect 8640 10580 8700 10600
rect 8770 10960 8830 10980
rect 8770 10600 8780 10960
rect 8820 10600 8830 10960
rect 8770 10580 8830 10600
rect 8900 10960 8960 10980
rect 8900 10600 8910 10960
rect 8950 10600 8960 10960
rect 8790 10520 8860 10540
rect 8790 10480 8810 10520
rect 8850 10480 8860 10520
rect 8790 10460 8860 10480
rect 8640 10410 8710 10430
rect 8900 10420 8960 10600
rect 9020 10770 9080 11040
rect 9730 11000 9810 11040
rect 9850 11000 9890 11040
rect 9930 11000 9970 11040
rect 10010 11000 10050 11040
rect 10090 11000 10130 11040
rect 10170 11000 10210 11040
rect 10250 11000 10290 11040
rect 10330 11000 10370 11040
rect 10410 11000 10450 11040
rect 10490 11000 10530 11040
rect 10570 11000 10610 11040
rect 10650 11000 10690 11040
rect 10730 11000 10770 11040
rect 10810 11000 10850 11040
rect 10890 11000 10930 11040
rect 10970 11000 11010 11040
rect 11050 11000 11090 11040
rect 11130 11000 11170 11040
rect 11210 11000 11250 11040
rect 11290 11000 11330 11040
rect 11370 11000 11410 11040
rect 11450 11000 11490 11040
rect 11530 11000 11570 11040
rect 11610 11000 11650 11040
rect 11690 11000 11730 11040
rect 11770 11000 11810 11040
rect 11850 11000 11890 11040
rect 11930 11000 11970 11040
rect 12010 11000 12050 11040
rect 12090 11000 12130 11040
rect 12170 11000 12210 11040
rect 12250 11000 12290 11040
rect 12330 11000 12370 11040
rect 12410 11000 12450 11040
rect 12490 11000 12530 11040
rect 12570 11000 12610 11040
rect 12650 11000 12690 11040
rect 12730 11000 12770 11040
rect 12810 11000 12850 11040
rect 12890 11000 12930 11040
rect 12970 11000 13010 11040
rect 13050 11000 13090 11040
rect 13130 11000 13170 11040
rect 13210 11000 13250 11040
rect 13290 11000 13330 11040
rect 13410 11000 13450 11040
rect 13490 11000 13530 11040
rect 13570 11000 13610 11040
rect 13650 11000 13690 11040
rect 13730 11000 13770 11040
rect 13810 11000 13850 11040
rect 13890 11000 13930 11040
rect 13970 11000 14010 11040
rect 14050 11000 14090 11040
rect 14130 11000 14170 11040
rect 14210 11000 14250 11040
rect 14290 11000 14330 11040
rect 14370 11000 14410 11040
rect 14450 11000 14490 11040
rect 14530 11000 14570 11040
rect 14610 11000 14650 11040
rect 14690 11000 14730 11040
rect 14770 11000 14810 11040
rect 14850 11000 14890 11040
rect 14930 11000 14970 11040
rect 15010 11000 15050 11040
rect 15090 11000 15130 11040
rect 15170 11000 15210 11040
rect 15250 11000 15290 11040
rect 15330 11000 15370 11040
rect 15410 11000 15450 11040
rect 15490 11000 15530 11040
rect 15570 11000 15610 11040
rect 15650 11000 15690 11040
rect 15730 11000 15770 11040
rect 15810 11000 15850 11040
rect 15890 11000 15930 11040
rect 15970 11000 16010 11040
rect 16050 11000 16090 11040
rect 16130 11000 16170 11040
rect 16210 11000 16250 11040
rect 16290 11000 16330 11040
rect 16370 11000 16410 11040
rect 16450 11000 16490 11040
rect 16530 11000 16570 11040
rect 16610 11000 16650 11040
rect 16690 11000 16730 11040
rect 16770 11000 16810 11040
rect 16850 11000 16890 11040
rect 16930 11000 16970 11040
rect 17010 11000 17050 11040
rect 17090 11000 17130 11040
rect 17170 11000 17210 11040
rect 17250 11000 17290 11040
rect 17330 11000 17370 11040
rect 17410 11000 17450 11040
rect 17490 11000 17530 11040
rect 17570 11000 17610 11040
rect 17650 11000 17690 11040
rect 17730 11000 17770 11040
rect 17810 11000 17850 11040
rect 17890 11000 17930 11040
rect 17970 11000 18010 11040
rect 18050 11000 18090 11040
rect 18130 11000 18170 11040
rect 18210 11000 18250 11040
rect 18290 11000 18330 11040
rect 18370 11000 18410 11040
rect 18450 11000 18490 11040
rect 18530 11000 18570 11040
rect 18610 11000 18650 11040
rect 18690 11000 18730 11040
rect 18770 11000 18810 11040
rect 18850 11000 18890 11040
rect 18930 11000 18970 11040
rect 19010 11000 19050 11040
rect 19090 11000 19130 11040
rect 19170 11000 19210 11040
rect 19250 11000 19290 11040
rect 19330 11000 19370 11040
rect 19410 11000 19450 11040
rect 19490 11000 19540 11040
rect 19580 11000 19620 11040
rect 19660 11000 19700 11040
rect 19740 11000 19780 11040
rect 19820 11000 19860 11040
rect 19900 11000 19940 11040
rect 19980 11000 20020 11040
rect 20060 11000 20110 11040
rect 20150 11000 20190 11040
rect 20230 11000 20270 11040
rect 20310 11000 20350 11040
rect 20390 11000 20430 11040
rect 20470 11000 20510 11040
rect 20550 11000 20590 11040
rect 20630 11000 20670 11040
rect 20710 11000 20750 11040
rect 20790 11000 20830 11040
rect 20870 11000 20910 11040
rect 20950 11000 20990 11040
rect 21030 11000 21070 11040
rect 21110 11000 21160 11040
rect 9730 10990 21160 11000
rect 9860 10910 9920 10990
rect 9020 10710 9590 10770
rect 9860 10750 9870 10910
rect 9910 10750 9920 10910
rect 9860 10730 9920 10750
rect 9970 10910 10030 10930
rect 9970 10750 9980 10910
rect 10020 10750 10030 10910
rect 9020 10650 9080 10710
rect 9020 10490 9030 10650
rect 9070 10490 9080 10650
rect 9020 10470 9080 10490
rect 9130 10650 9190 10670
rect 9130 10490 9140 10650
rect 9180 10490 9190 10650
rect 9130 10420 9190 10490
rect 9280 10650 9340 10710
rect 9280 10490 9290 10650
rect 9330 10490 9340 10650
rect 9280 10470 9340 10490
rect 9390 10650 9450 10670
rect 9390 10490 9400 10650
rect 9440 10490 9450 10650
rect 9390 10420 9450 10490
rect 9530 10650 9590 10710
rect 9840 10680 9930 10690
rect 9530 10490 9540 10650
rect 9580 10490 9590 10650
rect 9530 10470 9590 10490
rect 9640 10650 9700 10670
rect 9640 10490 9650 10650
rect 9690 10490 9700 10650
rect 9840 10640 9860 10680
rect 9900 10640 9930 10680
rect 9840 10630 9930 10640
rect 9640 10420 9700 10490
rect 8640 10370 8660 10410
rect 8700 10370 8710 10410
rect 8640 10350 8710 10370
rect 8770 10400 9090 10420
rect 8770 10360 8960 10400
rect 9000 10360 9040 10400
rect 9080 10360 9090 10400
rect 8770 10340 9090 10360
rect 9130 10400 9350 10420
rect 9130 10360 9160 10400
rect 9200 10360 9300 10400
rect 9340 10360 9350 10400
rect 9130 10340 9350 10360
rect 9390 10400 9600 10420
rect 9390 10360 9420 10400
rect 9460 10360 9550 10400
rect 9590 10360 9600 10400
rect 9390 10340 9600 10360
rect 9640 10400 9720 10420
rect 9640 10360 9670 10400
rect 9710 10360 9720 10400
rect 9640 10340 9720 10360
rect 9970 10390 10030 10750
rect 10080 10910 10140 10990
rect 10080 10750 10090 10910
rect 10130 10750 10140 10910
rect 10080 10730 10140 10750
rect 10510 10910 10570 10990
rect 10510 10550 10520 10910
rect 10560 10550 10570 10910
rect 10510 10530 10570 10550
rect 10770 10910 10830 10930
rect 10770 10550 10780 10910
rect 10820 10550 10830 10910
rect 11000 10910 11060 10990
rect 11000 10750 11010 10910
rect 11050 10750 11060 10910
rect 11000 10730 11060 10750
rect 11110 10910 11170 10930
rect 11110 10750 11120 10910
rect 11160 10750 11170 10910
rect 10670 10490 10730 10510
rect 10670 10450 10680 10490
rect 10720 10450 10730 10490
rect 10670 10430 10730 10450
rect 10410 10390 10470 10410
rect 10770 10390 10830 10550
rect 11110 10390 11170 10750
rect 11220 10910 11280 10990
rect 11220 10750 11230 10910
rect 11270 10750 11280 10910
rect 11220 10730 11280 10750
rect 11500 10910 11560 10990
rect 11500 10550 11510 10910
rect 11550 10550 11560 10910
rect 11500 10530 11560 10550
rect 11760 10910 11820 10930
rect 11760 10550 11770 10910
rect 11810 10550 11820 10910
rect 11990 10910 12050 10990
rect 11990 10750 12000 10910
rect 12040 10750 12050 10910
rect 11990 10730 12050 10750
rect 12100 10910 12160 10930
rect 12100 10750 12110 10910
rect 12150 10750 12160 10910
rect 11660 10490 11720 10510
rect 11660 10450 11670 10490
rect 11710 10450 11720 10490
rect 11660 10430 11720 10450
rect 11400 10390 11460 10410
rect 11760 10390 11820 10550
rect 12100 10390 12160 10750
rect 12210 10910 12270 10990
rect 12210 10750 12220 10910
rect 12260 10750 12270 10910
rect 12210 10730 12270 10750
rect 12500 10910 12560 10990
rect 12500 10550 12510 10910
rect 12550 10550 12560 10910
rect 12500 10530 12560 10550
rect 12760 10910 12820 10930
rect 12760 10550 12770 10910
rect 12810 10550 12820 10910
rect 12990 10910 13050 10990
rect 12990 10750 13000 10910
rect 13040 10750 13050 10910
rect 12990 10730 13050 10750
rect 13100 10910 13160 10930
rect 13100 10750 13110 10910
rect 13150 10750 13160 10910
rect 12660 10490 12720 10510
rect 12660 10450 12670 10490
rect 12710 10450 12720 10490
rect 12660 10430 12720 10450
rect 12400 10390 12460 10410
rect 12760 10390 12820 10550
rect 13100 10410 13160 10750
rect 13210 10910 13270 10990
rect 13210 10750 13220 10910
rect 13260 10750 13270 10910
rect 13210 10730 13270 10750
rect 13330 10630 13390 10990
rect 13330 10470 13340 10630
rect 13380 10470 13390 10630
rect 13330 10450 13390 10470
rect 13440 10630 13500 10650
rect 13440 10470 13450 10630
rect 13490 10470 13500 10630
rect 13100 10390 13400 10410
rect 9970 10380 10220 10390
rect 9970 10340 10160 10380
rect 10200 10340 10220 10380
rect 8220 9720 8280 9740
rect 8640 10280 8700 10300
rect 8640 9820 8650 10280
rect 8690 9820 8700 10280
rect 8640 9730 8700 9820
rect 8770 10280 8830 10340
rect 8770 9820 8780 10280
rect 8820 9820 8830 10280
rect 8770 9800 8830 9820
rect 8900 10280 8960 10300
rect 8900 9820 8910 10280
rect 8950 9820 8960 10280
rect 8900 9730 8960 9820
rect 9020 10280 9080 10300
rect 9020 9820 9030 10280
rect 9070 9820 9080 10280
rect 9020 9730 9080 9820
rect 9130 10280 9190 10340
rect 9130 9820 9140 10280
rect 9180 9820 9190 10280
rect 9130 9800 9190 9820
rect 9280 10280 9340 10300
rect 9280 9820 9290 10280
rect 9330 9820 9340 10280
rect 9280 9730 9340 9820
rect 9390 10280 9450 10340
rect 9390 9820 9400 10280
rect 9440 9820 9450 10280
rect 9390 9800 9450 9820
rect 9530 10280 9590 10300
rect 9530 9820 9540 10280
rect 9580 9820 9590 10280
rect 9530 9730 9590 9820
rect 9640 10280 9700 10340
rect 9970 10330 10220 10340
rect 10410 10350 10420 10390
rect 10460 10350 10470 10390
rect 10410 10330 10470 10350
rect 10640 10380 11070 10390
rect 10640 10340 10920 10380
rect 10960 10340 11000 10380
rect 11040 10340 11070 10380
rect 10640 10330 11070 10340
rect 11110 10380 11350 10390
rect 11110 10340 11300 10380
rect 11340 10340 11350 10380
rect 11110 10330 11350 10340
rect 11400 10350 11410 10390
rect 11450 10350 11460 10390
rect 11400 10330 11460 10350
rect 11630 10380 12060 10390
rect 11630 10340 11910 10380
rect 11950 10340 11990 10380
rect 12030 10340 12060 10380
rect 11630 10330 12060 10340
rect 12100 10380 12340 10390
rect 12100 10340 12290 10380
rect 12330 10340 12340 10380
rect 12100 10330 12340 10340
rect 12400 10350 12410 10390
rect 12450 10350 12460 10390
rect 12400 10330 12460 10350
rect 12630 10380 13060 10390
rect 12630 10340 12910 10380
rect 12950 10340 12990 10380
rect 13030 10340 13060 10380
rect 12630 10330 13060 10340
rect 13100 10350 13270 10390
rect 13310 10350 13350 10390
rect 13390 10350 13400 10390
rect 13100 10330 13400 10350
rect 13440 10390 13500 10470
rect 13560 10630 13620 10650
rect 13560 10470 13570 10630
rect 13610 10470 13620 10630
rect 13560 10450 13620 10470
rect 13670 10630 13730 10990
rect 13670 10470 13680 10630
rect 13720 10470 13730 10630
rect 13670 10450 13730 10470
rect 13780 10630 13840 10650
rect 13780 10470 13790 10630
rect 13830 10470 13840 10630
rect 13440 10350 13450 10390
rect 13490 10350 13500 10390
rect 9640 9820 9650 10280
rect 9690 9820 9700 10280
rect 9640 9800 9700 9820
rect 9860 10270 9920 10290
rect 9860 9810 9870 10270
rect 9910 9810 9920 10270
rect 9860 9730 9920 9810
rect 9970 10270 10030 10330
rect 9970 9810 9980 10270
rect 10020 9810 10030 10270
rect 9970 9790 10030 9810
rect 10080 10270 10140 10290
rect 10080 9810 10090 10270
rect 10130 9810 10140 10270
rect 10080 9730 10140 9810
rect 10510 10270 10570 10290
rect 10510 9810 10520 10270
rect 10560 9810 10570 10270
rect 10510 9730 10570 9810
rect 10640 10270 10700 10330
rect 10640 9810 10650 10270
rect 10690 9810 10700 10270
rect 10640 9790 10700 9810
rect 10770 10270 10830 10290
rect 10770 9810 10780 10270
rect 10820 9810 10830 10270
rect 10770 9730 10830 9810
rect 11000 10270 11060 10290
rect 11000 9810 11010 10270
rect 11050 9810 11060 10270
rect 11000 9730 11060 9810
rect 11110 10270 11170 10330
rect 11110 9810 11120 10270
rect 11160 9810 11170 10270
rect 11110 9790 11170 9810
rect 11220 10270 11280 10290
rect 11220 9810 11230 10270
rect 11270 9810 11280 10270
rect 11220 9730 11280 9810
rect 11500 10270 11560 10290
rect 11500 9810 11510 10270
rect 11550 9810 11560 10270
rect 11500 9730 11560 9810
rect 11630 10270 11690 10330
rect 11630 9810 11640 10270
rect 11680 9810 11690 10270
rect 11630 9790 11690 9810
rect 11760 10270 11820 10290
rect 11760 9810 11770 10270
rect 11810 9810 11820 10270
rect 11760 9730 11820 9810
rect 11990 10270 12050 10290
rect 11990 9810 12000 10270
rect 12040 9810 12050 10270
rect 11990 9730 12050 9810
rect 12100 10270 12160 10330
rect 12100 9810 12110 10270
rect 12150 9810 12160 10270
rect 12100 9790 12160 9810
rect 12210 10270 12270 10290
rect 12210 9810 12220 10270
rect 12260 9810 12270 10270
rect 12210 9730 12270 9810
rect 12500 10270 12560 10290
rect 12500 9810 12510 10270
rect 12550 9810 12560 10270
rect 12500 9730 12560 9810
rect 12630 10270 12690 10330
rect 12630 9810 12640 10270
rect 12680 9810 12690 10270
rect 12630 9790 12690 9810
rect 12760 10270 12820 10290
rect 12760 9810 12770 10270
rect 12810 9810 12820 10270
rect 12760 9730 12820 9810
rect 12990 10270 13050 10290
rect 12990 9810 13000 10270
rect 13040 9810 13050 10270
rect 12990 9730 13050 9810
rect 13100 10270 13160 10330
rect 13100 9810 13110 10270
rect 13150 9810 13160 10270
rect 13100 9790 13160 9810
rect 13210 10270 13270 10290
rect 13210 9810 13220 10270
rect 13260 9810 13270 10270
rect 13210 9730 13270 9810
rect 13330 10270 13390 10290
rect 13330 9810 13340 10270
rect 13380 9810 13390 10270
rect 13330 9730 13390 9810
rect 13440 10270 13500 10350
rect 13570 10390 13630 10410
rect 13570 10350 13580 10390
rect 13620 10350 13630 10390
rect 13570 10330 13630 10350
rect 13780 10390 13840 10470
rect 13900 10630 13960 10650
rect 13900 10470 13910 10630
rect 13950 10470 13960 10630
rect 13900 10450 13960 10470
rect 14010 10630 14070 10990
rect 14010 10470 14020 10630
rect 14060 10470 14070 10630
rect 14010 10450 14070 10470
rect 14120 10630 14180 10650
rect 14120 10470 14130 10630
rect 14170 10470 14180 10630
rect 14120 10450 14180 10470
rect 14230 10630 14290 10990
rect 14230 10470 14240 10630
rect 14280 10470 14290 10630
rect 14230 10450 14290 10470
rect 14340 10630 14400 10650
rect 14340 10470 14350 10630
rect 14390 10470 14400 10630
rect 13780 10350 13790 10390
rect 13830 10350 13840 10390
rect 13440 9810 13450 10270
rect 13490 9810 13500 10270
rect 13440 9790 13500 9810
rect 13560 10270 13620 10290
rect 13560 9810 13570 10270
rect 13610 9810 13620 10270
rect 13560 9790 13620 9810
rect 13670 10270 13730 10290
rect 13670 9810 13680 10270
rect 13720 9810 13730 10270
rect 13670 9730 13730 9810
rect 13780 10270 13840 10350
rect 13910 10390 13970 10410
rect 13910 10350 13920 10390
rect 13960 10350 13970 10390
rect 13910 10330 13970 10350
rect 14340 10390 14400 10470
rect 14460 10630 14520 10650
rect 14460 10470 14470 10630
rect 14510 10470 14520 10630
rect 14460 10450 14520 10470
rect 14570 10630 14630 10990
rect 14570 10470 14580 10630
rect 14620 10470 14630 10630
rect 14570 10450 14630 10470
rect 14680 10630 14740 10650
rect 14680 10470 14690 10630
rect 14730 10470 14740 10630
rect 14680 10450 14740 10470
rect 14790 10630 14850 10990
rect 14790 10470 14800 10630
rect 14840 10470 14850 10630
rect 14790 10450 14850 10470
rect 14900 10630 14960 10650
rect 14900 10470 14910 10630
rect 14950 10470 14960 10630
rect 14900 10450 14960 10470
rect 15010 10630 15070 10990
rect 15010 10470 15020 10630
rect 15060 10470 15070 10630
rect 15010 10450 15070 10470
rect 15120 10630 15180 10650
rect 15120 10470 15130 10630
rect 15170 10470 15180 10630
rect 15120 10450 15180 10470
rect 15230 10630 15290 10990
rect 15230 10470 15240 10630
rect 15280 10470 15290 10630
rect 15230 10450 15290 10470
rect 15340 10630 15400 10650
rect 15340 10470 15350 10630
rect 15390 10470 15400 10630
rect 14340 10350 14350 10390
rect 14390 10350 14400 10390
rect 13780 9810 13790 10270
rect 13830 9810 13840 10270
rect 13780 9790 13840 9810
rect 13900 10270 13960 10290
rect 13900 9810 13910 10270
rect 13950 9810 13960 10270
rect 13900 9790 13960 9810
rect 14010 10270 14070 10290
rect 14010 9810 14020 10270
rect 14060 9810 14070 10270
rect 14010 9730 14070 9810
rect 14120 10270 14180 10290
rect 14120 9810 14130 10270
rect 14170 9810 14180 10270
rect 14120 9790 14180 9810
rect 14230 10270 14290 10290
rect 14230 9810 14240 10270
rect 14280 9810 14290 10270
rect 14230 9730 14290 9810
rect 14340 10270 14400 10350
rect 14470 10390 14530 10410
rect 14470 10350 14480 10390
rect 14520 10350 14530 10390
rect 14470 10330 14530 10350
rect 15340 10390 15400 10470
rect 15520 10630 15580 10650
rect 15520 10470 15530 10630
rect 15570 10470 15580 10630
rect 15520 10450 15580 10470
rect 15630 10630 15690 10990
rect 15630 10470 15640 10630
rect 15680 10470 15690 10630
rect 15630 10450 15690 10470
rect 15740 10630 15800 10650
rect 15740 10470 15750 10630
rect 15790 10470 15800 10630
rect 15740 10450 15800 10470
rect 15850 10630 15910 10990
rect 15850 10470 15860 10630
rect 15900 10470 15910 10630
rect 15850 10450 15910 10470
rect 15960 10630 16020 10650
rect 15960 10470 15970 10630
rect 16010 10470 16020 10630
rect 15960 10450 16020 10470
rect 16070 10630 16130 10990
rect 16070 10470 16080 10630
rect 16120 10470 16130 10630
rect 16070 10450 16130 10470
rect 16180 10630 16240 10650
rect 16180 10470 16190 10630
rect 16230 10470 16240 10630
rect 16180 10450 16240 10470
rect 16290 10630 16350 10990
rect 16290 10470 16300 10630
rect 16340 10470 16350 10630
rect 16290 10450 16350 10470
rect 16400 10630 16460 10650
rect 16400 10470 16410 10630
rect 16450 10470 16460 10630
rect 16400 10450 16460 10470
rect 16510 10630 16570 10990
rect 16510 10470 16520 10630
rect 16560 10470 16570 10630
rect 16510 10450 16570 10470
rect 16620 10630 16680 10650
rect 16620 10470 16630 10630
rect 16670 10470 16680 10630
rect 16620 10450 16680 10470
rect 16730 10630 16790 10990
rect 16730 10470 16740 10630
rect 16780 10470 16790 10630
rect 16730 10450 16790 10470
rect 16840 10630 16900 10650
rect 16840 10470 16850 10630
rect 16890 10470 16900 10630
rect 16840 10450 16900 10470
rect 16950 10630 17010 10990
rect 16950 10470 16960 10630
rect 17000 10470 17010 10630
rect 16950 10450 17010 10470
rect 17060 10630 17120 10650
rect 17060 10470 17070 10630
rect 17110 10470 17120 10630
rect 17060 10450 17120 10470
rect 17170 10630 17230 10990
rect 17170 10470 17180 10630
rect 17220 10470 17230 10630
rect 17170 10450 17230 10470
rect 17280 10630 17340 10650
rect 17280 10470 17290 10630
rect 17330 10470 17340 10630
rect 17280 10410 17340 10470
rect 17470 10630 17530 10650
rect 17470 10470 17480 10630
rect 17520 10470 17530 10630
rect 17470 10450 17530 10470
rect 17580 10630 17640 10990
rect 17580 10470 17590 10630
rect 17630 10470 17640 10630
rect 17580 10450 17640 10470
rect 17690 10630 17750 10650
rect 17690 10470 17700 10630
rect 17740 10470 17750 10630
rect 17690 10450 17750 10470
rect 17800 10630 17860 10990
rect 17800 10470 17810 10630
rect 17850 10470 17860 10630
rect 17800 10450 17860 10470
rect 17910 10630 17970 10650
rect 17910 10470 17920 10630
rect 17960 10470 17970 10630
rect 17910 10450 17970 10470
rect 18020 10630 18080 10990
rect 18020 10470 18030 10630
rect 18070 10470 18080 10630
rect 18020 10450 18080 10470
rect 18130 10630 18190 10650
rect 18130 10470 18140 10630
rect 18180 10470 18190 10630
rect 18130 10450 18190 10470
rect 18240 10630 18300 10990
rect 18240 10470 18250 10630
rect 18290 10470 18300 10630
rect 18240 10450 18300 10470
rect 18350 10630 18410 10650
rect 18350 10470 18360 10630
rect 18400 10470 18410 10630
rect 18350 10450 18410 10470
rect 18460 10630 18520 10990
rect 18460 10470 18470 10630
rect 18510 10470 18520 10630
rect 18460 10450 18520 10470
rect 18570 10630 18630 10650
rect 18570 10470 18580 10630
rect 18620 10470 18630 10630
rect 18570 10450 18630 10470
rect 18680 10630 18740 10990
rect 18680 10470 18690 10630
rect 18730 10470 18740 10630
rect 18680 10450 18740 10470
rect 18790 10630 18850 10650
rect 18790 10470 18800 10630
rect 18840 10470 18850 10630
rect 18790 10450 18850 10470
rect 18900 10630 18960 10990
rect 18900 10470 18910 10630
rect 18950 10470 18960 10630
rect 18900 10450 18960 10470
rect 19010 10630 19070 10650
rect 19010 10470 19020 10630
rect 19060 10470 19070 10630
rect 19010 10450 19070 10470
rect 19120 10630 19180 10990
rect 19120 10470 19130 10630
rect 19170 10470 19180 10630
rect 19120 10450 19180 10470
rect 19230 10630 19290 10650
rect 19230 10470 19240 10630
rect 19280 10470 19290 10630
rect 19230 10450 19290 10470
rect 19340 10630 19400 10990
rect 19340 10470 19350 10630
rect 19390 10470 19400 10630
rect 19340 10450 19400 10470
rect 19450 10630 19510 10650
rect 19450 10470 19460 10630
rect 19500 10470 19510 10630
rect 19450 10450 19510 10470
rect 19560 10630 19620 10990
rect 19560 10470 19570 10630
rect 19610 10470 19620 10630
rect 19560 10450 19620 10470
rect 19670 10630 19730 10650
rect 19670 10470 19680 10630
rect 19720 10470 19730 10630
rect 19670 10450 19730 10470
rect 19780 10630 19840 10990
rect 19780 10470 19790 10630
rect 19830 10470 19840 10630
rect 19780 10450 19840 10470
rect 19890 10630 19950 10650
rect 19890 10470 19900 10630
rect 19940 10470 19950 10630
rect 19890 10450 19950 10470
rect 20000 10630 20060 10990
rect 20000 10470 20010 10630
rect 20050 10470 20060 10630
rect 20000 10450 20060 10470
rect 20110 10630 20170 10650
rect 20110 10470 20120 10630
rect 20160 10470 20170 10630
rect 20110 10450 20170 10470
rect 20220 10630 20280 10990
rect 20220 10470 20230 10630
rect 20270 10470 20280 10630
rect 20220 10450 20280 10470
rect 20330 10630 20390 10650
rect 20330 10470 20340 10630
rect 20380 10470 20390 10630
rect 20330 10450 20390 10470
rect 20440 10630 20500 10990
rect 20440 10470 20450 10630
rect 20490 10470 20500 10630
rect 20440 10450 20500 10470
rect 20550 10630 20610 10650
rect 20550 10470 20560 10630
rect 20600 10470 20610 10630
rect 20550 10450 20610 10470
rect 20660 10630 20720 10990
rect 20660 10470 20670 10630
rect 20710 10470 20720 10630
rect 20660 10450 20720 10470
rect 20770 10630 20830 10650
rect 20770 10470 20780 10630
rect 20820 10470 20830 10630
rect 20770 10450 20830 10470
rect 20880 10630 20940 10990
rect 20880 10470 20890 10630
rect 20930 10470 20940 10630
rect 20880 10450 20940 10470
rect 20990 10630 21050 10650
rect 20990 10470 21000 10630
rect 21040 10470 21050 10630
rect 20990 10410 21050 10470
rect 15340 10350 15350 10390
rect 15390 10350 15400 10390
rect 14340 9810 14350 10270
rect 14390 9810 14400 10270
rect 14340 9790 14400 9810
rect 14460 10270 14520 10290
rect 14460 9810 14470 10270
rect 14510 9810 14520 10270
rect 14460 9790 14520 9810
rect 14570 10270 14630 10290
rect 14570 9810 14580 10270
rect 14620 9810 14630 10270
rect 14570 9730 14630 9810
rect 14680 10270 14740 10290
rect 14680 9810 14690 10270
rect 14730 9810 14740 10270
rect 14680 9790 14740 9810
rect 14790 10270 14850 10290
rect 14790 9810 14800 10270
rect 14840 9810 14850 10270
rect 14790 9730 14850 9810
rect 14900 10270 14960 10290
rect 14900 9810 14910 10270
rect 14950 9810 14960 10270
rect 14900 9790 14960 9810
rect 15010 10270 15070 10290
rect 15010 9810 15020 10270
rect 15060 9810 15070 10270
rect 15010 9730 15070 9810
rect 15120 10270 15180 10290
rect 15120 9810 15130 10270
rect 15170 9810 15180 10270
rect 15120 9790 15180 9810
rect 15230 10270 15290 10290
rect 15230 9810 15240 10270
rect 15280 9810 15290 10270
rect 15230 9730 15290 9810
rect 15340 10270 15400 10350
rect 15530 10390 15590 10410
rect 15530 10350 15540 10390
rect 15580 10350 15590 10390
rect 15530 10330 15590 10350
rect 17280 10400 17410 10410
rect 17280 10350 17340 10400
rect 17390 10350 17410 10400
rect 17280 10340 17410 10350
rect 17470 10390 17540 10410
rect 17470 10350 17490 10390
rect 17530 10350 17540 10390
rect 15340 9810 15350 10270
rect 15390 9810 15400 10270
rect 15340 9790 15400 9810
rect 15520 10270 15580 10290
rect 15520 9810 15530 10270
rect 15570 9810 15580 10270
rect 15520 9790 15580 9810
rect 15630 10270 15690 10290
rect 15630 9810 15640 10270
rect 15680 9810 15690 10270
rect 15630 9730 15690 9810
rect 15740 10270 15800 10290
rect 15740 9810 15750 10270
rect 15790 9810 15800 10270
rect 15740 9790 15800 9810
rect 15850 10270 15910 10290
rect 15850 9810 15860 10270
rect 15900 9810 15910 10270
rect 15850 9730 15910 9810
rect 15960 10270 16020 10290
rect 15960 9810 15970 10270
rect 16010 9810 16020 10270
rect 15960 9790 16020 9810
rect 16070 10270 16130 10290
rect 16070 9810 16080 10270
rect 16120 9810 16130 10270
rect 16070 9730 16130 9810
rect 16180 10270 16240 10290
rect 16180 9810 16190 10270
rect 16230 9810 16240 10270
rect 16180 9790 16240 9810
rect 16290 10270 16350 10290
rect 16290 9810 16300 10270
rect 16340 9810 16350 10270
rect 16290 9730 16350 9810
rect 16400 10270 16460 10290
rect 16400 9810 16410 10270
rect 16450 9810 16460 10270
rect 16400 9790 16460 9810
rect 16510 10270 16570 10290
rect 16510 9810 16520 10270
rect 16560 9810 16570 10270
rect 16510 9730 16570 9810
rect 16620 10270 16680 10290
rect 16620 9810 16630 10270
rect 16670 9810 16680 10270
rect 16620 9790 16680 9810
rect 16730 10270 16790 10290
rect 16730 9810 16740 10270
rect 16780 9810 16790 10270
rect 16730 9730 16790 9810
rect 16840 10270 16900 10290
rect 16840 9810 16850 10270
rect 16890 9810 16900 10270
rect 16840 9790 16900 9810
rect 16950 10270 17010 10290
rect 16950 9810 16960 10270
rect 17000 9810 17010 10270
rect 16950 9730 17010 9810
rect 17060 10270 17120 10290
rect 17060 9810 17070 10270
rect 17110 9810 17120 10270
rect 17060 9790 17120 9810
rect 17170 10270 17230 10290
rect 17170 9810 17180 10270
rect 17220 9810 17230 10270
rect 17170 9730 17230 9810
rect 17280 10270 17340 10340
rect 17470 10330 17540 10350
rect 20990 10400 21120 10410
rect 20990 10350 21050 10400
rect 21100 10350 21120 10400
rect 20990 10340 21120 10350
rect 17280 9810 17290 10270
rect 17330 9810 17340 10270
rect 17280 9790 17340 9810
rect 17470 10270 17530 10290
rect 17470 9810 17480 10270
rect 17520 9810 17530 10270
rect 17470 9790 17530 9810
rect 17580 10270 17640 10290
rect 17580 9810 17590 10270
rect 17630 9810 17640 10270
rect 17580 9730 17640 9810
rect 17690 10270 17750 10290
rect 17690 9810 17700 10270
rect 17740 9810 17750 10270
rect 17690 9790 17750 9810
rect 17800 10270 17860 10290
rect 17800 9810 17810 10270
rect 17850 9810 17860 10270
rect 17800 9730 17860 9810
rect 17910 10270 17970 10290
rect 17910 9810 17920 10270
rect 17960 9810 17970 10270
rect 17910 9790 17970 9810
rect 18020 10270 18080 10290
rect 18020 9810 18030 10270
rect 18070 9810 18080 10270
rect 18020 9730 18080 9810
rect 18130 10270 18190 10290
rect 18130 9810 18140 10270
rect 18180 9810 18190 10270
rect 18130 9790 18190 9810
rect 18240 10270 18300 10290
rect 18240 9810 18250 10270
rect 18290 9810 18300 10270
rect 18240 9730 18300 9810
rect 18350 10270 18410 10290
rect 18350 9810 18360 10270
rect 18400 9810 18410 10270
rect 18350 9790 18410 9810
rect 18460 10270 18520 10290
rect 18460 9810 18470 10270
rect 18510 9810 18520 10270
rect 18460 9730 18520 9810
rect 18570 10270 18630 10290
rect 18570 9810 18580 10270
rect 18620 9810 18630 10270
rect 18570 9790 18630 9810
rect 18680 10270 18740 10290
rect 18680 9810 18690 10270
rect 18730 9810 18740 10270
rect 18680 9730 18740 9810
rect 18790 10270 18850 10290
rect 18790 9810 18800 10270
rect 18840 9810 18850 10270
rect 18790 9790 18850 9810
rect 18900 10270 18960 10290
rect 18900 9810 18910 10270
rect 18950 9810 18960 10270
rect 18900 9730 18960 9810
rect 19010 10270 19070 10290
rect 19010 9810 19020 10270
rect 19060 9810 19070 10270
rect 19010 9790 19070 9810
rect 19120 10270 19180 10290
rect 19120 9810 19130 10270
rect 19170 9810 19180 10270
rect 19120 9730 19180 9810
rect 19230 10270 19290 10290
rect 19230 9810 19240 10270
rect 19280 9810 19290 10270
rect 19230 9790 19290 9810
rect 19340 10270 19400 10290
rect 19340 9810 19350 10270
rect 19390 9810 19400 10270
rect 19340 9730 19400 9810
rect 19450 10270 19510 10290
rect 19450 9810 19460 10270
rect 19500 9810 19510 10270
rect 19450 9790 19510 9810
rect 19560 10270 19620 10290
rect 19560 9810 19570 10270
rect 19610 9810 19620 10270
rect 19560 9730 19620 9810
rect 19670 10270 19730 10290
rect 19670 9810 19680 10270
rect 19720 9810 19730 10270
rect 19670 9790 19730 9810
rect 19780 10270 19840 10290
rect 19780 9810 19790 10270
rect 19830 9810 19840 10270
rect 19780 9730 19840 9810
rect 19890 10270 19950 10290
rect 19890 9810 19900 10270
rect 19940 9810 19950 10270
rect 19890 9790 19950 9810
rect 20000 10270 20060 10290
rect 20000 9810 20010 10270
rect 20050 9810 20060 10270
rect 20000 9730 20060 9810
rect 20110 10270 20170 10290
rect 20110 9810 20120 10270
rect 20160 9810 20170 10270
rect 20110 9790 20170 9810
rect 20220 10270 20280 10290
rect 20220 9810 20230 10270
rect 20270 9810 20280 10270
rect 20220 9730 20280 9810
rect 20330 10270 20390 10290
rect 20330 9810 20340 10270
rect 20380 9810 20390 10270
rect 20330 9790 20390 9810
rect 20440 10270 20500 10290
rect 20440 9810 20450 10270
rect 20490 9810 20500 10270
rect 20440 9730 20500 9810
rect 20550 10270 20610 10290
rect 20550 9810 20560 10270
rect 20600 9810 20610 10270
rect 20550 9790 20610 9810
rect 20660 10270 20720 10290
rect 20660 9810 20670 10270
rect 20710 9810 20720 10270
rect 20660 9730 20720 9810
rect 20770 10270 20830 10290
rect 20770 9810 20780 10270
rect 20820 9810 20830 10270
rect 20770 9790 20830 9810
rect 20880 10270 20940 10290
rect 20880 9810 20890 10270
rect 20930 9810 20940 10270
rect 20880 9730 20940 9810
rect 20990 10270 21050 10340
rect 20990 9810 21000 10270
rect 21040 9810 21050 10270
rect 20990 9790 21050 9810
rect 8470 9720 21120 9730
rect 8470 9680 8520 9720
rect 8560 9680 8600 9720
rect 8640 9680 8680 9720
rect 8720 9680 8760 9720
rect 8800 9680 8840 9720
rect 8880 9680 8920 9720
rect 8960 9680 9000 9720
rect 9040 9680 9080 9720
rect 9120 9680 9160 9720
rect 9200 9680 9240 9720
rect 9280 9680 9320 9720
rect 9360 9680 9400 9720
rect 9440 9680 9480 9720
rect 9520 9680 9560 9720
rect 9600 9680 9640 9720
rect 9680 9680 9720 9720
rect 9760 9680 9800 9720
rect 9840 9680 9890 9720
rect 9930 9680 9970 9720
rect 10010 9680 10050 9720
rect 10090 9680 10130 9720
rect 10170 9680 10210 9720
rect 10250 9680 10290 9720
rect 10330 9680 10370 9720
rect 10410 9680 10450 9720
rect 10490 9680 10530 9720
rect 10570 9680 10610 9720
rect 10650 9680 10690 9720
rect 10730 9680 10770 9720
rect 10810 9680 10850 9720
rect 10890 9680 10930 9720
rect 10970 9680 11010 9720
rect 11050 9680 11090 9720
rect 11130 9680 11170 9720
rect 11210 9680 11250 9720
rect 11290 9680 11330 9720
rect 11370 9680 11410 9720
rect 11450 9680 11490 9720
rect 11530 9680 11570 9720
rect 11610 9680 11650 9720
rect 11690 9680 11730 9720
rect 11770 9680 11810 9720
rect 11850 9680 11890 9720
rect 11930 9680 11970 9720
rect 12010 9680 12050 9720
rect 12090 9680 12130 9720
rect 12170 9680 12210 9720
rect 12250 9680 12290 9720
rect 12330 9680 12370 9720
rect 12410 9680 12450 9720
rect 12490 9680 12530 9720
rect 12570 9680 12610 9720
rect 12650 9680 12690 9720
rect 12730 9680 12770 9720
rect 12810 9680 12850 9720
rect 12890 9680 12930 9720
rect 12970 9680 13010 9720
rect 13050 9680 13090 9720
rect 13130 9680 13170 9720
rect 13210 9680 13250 9720
rect 13290 9680 13330 9720
rect 13370 9680 13410 9720
rect 13450 9680 13490 9720
rect 13530 9680 13570 9720
rect 13610 9680 13650 9720
rect 13690 9680 13730 9720
rect 13770 9680 13810 9720
rect 13850 9680 13890 9720
rect 13930 9680 13970 9720
rect 14010 9680 14050 9720
rect 14090 9680 14130 9720
rect 14170 9680 14210 9720
rect 14250 9680 14290 9720
rect 14330 9680 14370 9720
rect 14410 9680 14450 9720
rect 14490 9680 14530 9720
rect 14570 9680 14610 9720
rect 14650 9680 14690 9720
rect 14730 9680 14770 9720
rect 14810 9680 14850 9720
rect 14890 9680 14930 9720
rect 14970 9680 15010 9720
rect 15050 9680 15090 9720
rect 15130 9680 15170 9720
rect 15210 9680 15250 9720
rect 15290 9680 15330 9720
rect 15370 9680 15410 9720
rect 15450 9680 15490 9720
rect 15530 9680 15570 9720
rect 15610 9680 15650 9720
rect 15690 9680 15730 9720
rect 15770 9680 15810 9720
rect 15850 9680 15890 9720
rect 15930 9680 15970 9720
rect 16010 9680 16050 9720
rect 16090 9680 16130 9720
rect 16170 9680 16210 9720
rect 16250 9680 16290 9720
rect 16330 9680 16370 9720
rect 16410 9680 16450 9720
rect 16490 9680 16530 9720
rect 16570 9680 16610 9720
rect 16650 9680 16690 9720
rect 16730 9680 16770 9720
rect 16810 9680 16850 9720
rect 16890 9680 16930 9720
rect 16970 9680 17010 9720
rect 17050 9680 17090 9720
rect 17130 9680 17170 9720
rect 17210 9680 17250 9720
rect 17290 9680 17330 9720
rect 17370 9680 17410 9720
rect 17450 9680 17490 9720
rect 17530 9680 17570 9720
rect 17610 9680 17650 9720
rect 17690 9680 17730 9720
rect 17770 9680 17810 9720
rect 17850 9680 17890 9720
rect 17930 9680 17970 9720
rect 18010 9680 18050 9720
rect 18090 9680 18130 9720
rect 18170 9680 18210 9720
rect 18250 9680 18290 9720
rect 18330 9680 18370 9720
rect 18410 9680 18450 9720
rect 18490 9680 18530 9720
rect 18570 9680 18610 9720
rect 18650 9680 18690 9720
rect 18730 9680 18770 9720
rect 18810 9680 18850 9720
rect 18890 9680 18930 9720
rect 18970 9680 19010 9720
rect 19050 9680 19090 9720
rect 19130 9680 19170 9720
rect 19210 9680 19250 9720
rect 19290 9680 19330 9720
rect 19370 9680 19410 9720
rect 19450 9680 19490 9720
rect 19530 9680 19570 9720
rect 19610 9680 19650 9720
rect 19690 9680 19730 9720
rect 19770 9680 19810 9720
rect 19850 9680 19890 9720
rect 19930 9680 19970 9720
rect 20010 9680 20050 9720
rect 20090 9680 20130 9720
rect 20170 9680 20210 9720
rect 20250 9680 20290 9720
rect 20330 9680 20370 9720
rect 20410 9680 20450 9720
rect 20490 9680 20530 9720
rect 20570 9680 20610 9720
rect 20650 9680 20690 9720
rect 20730 9680 20770 9720
rect 20810 9680 20850 9720
rect 20890 9680 20930 9720
rect 20970 9680 21010 9720
rect 21050 9680 21120 9720
rect 8470 9670 21120 9680
rect 8470 9650 8530 9670
rect 7710 9630 8530 9650
rect 7710 9590 7740 9630
rect 7780 9590 7820 9630
rect 7860 9590 7900 9630
rect 7940 9590 7980 9630
rect 8020 9590 8060 9630
rect 8100 9590 8140 9630
rect 8180 9590 8220 9630
rect 8260 9590 8300 9630
rect 8340 9590 8380 9630
rect 8420 9590 8460 9630
rect 8500 9590 8530 9630
rect 7710 9570 8530 9590
rect 13190 8630 13300 8640
rect 13190 8580 13220 8630
rect 13270 8580 13300 8630
rect 13190 8570 13300 8580
rect 13390 8490 13600 8510
rect 13390 8480 13430 8490
rect 9890 8430 13430 8480
rect 9900 8240 9960 8260
rect 9900 7080 9910 8240
rect 9950 7080 9960 8240
rect 9900 6990 9960 7080
rect 10010 8240 10070 8430
rect 10010 7080 10020 8240
rect 10060 7080 10070 8240
rect 10010 7060 10070 7080
rect 10120 8240 10180 8260
rect 10120 7080 10130 8240
rect 10170 7080 10180 8240
rect 10120 6990 10180 7080
rect 10230 8240 10290 8430
rect 10230 7080 10240 8240
rect 10280 7080 10290 8240
rect 10230 7060 10290 7080
rect 10340 8240 10400 8260
rect 10340 7080 10350 8240
rect 10390 7080 10400 8240
rect 10340 6990 10400 7080
rect 10450 8240 10510 8430
rect 10450 7080 10460 8240
rect 10500 7080 10510 8240
rect 10450 7060 10510 7080
rect 10560 8240 10620 8260
rect 10560 7080 10570 8240
rect 10610 7080 10620 8240
rect 10560 6990 10620 7080
rect 10670 8240 10730 8430
rect 10670 7080 10680 8240
rect 10720 7080 10730 8240
rect 10670 7060 10730 7080
rect 10780 8240 10840 8260
rect 10780 7080 10790 8240
rect 10830 7080 10840 8240
rect 10780 6990 10840 7080
rect 10890 8240 10950 8430
rect 10890 7080 10900 8240
rect 10940 7080 10950 8240
rect 10890 7060 10950 7080
rect 11000 8240 11060 8260
rect 11000 7080 11010 8240
rect 11050 7080 11060 8240
rect 11000 6990 11060 7080
rect 11110 8240 11170 8430
rect 11110 7080 11120 8240
rect 11160 7080 11170 8240
rect 11110 7060 11170 7080
rect 11220 8240 11280 8260
rect 11220 7080 11230 8240
rect 11270 7080 11280 8240
rect 11220 6990 11280 7080
rect 11330 8240 11390 8430
rect 11330 7080 11340 8240
rect 11380 7080 11390 8240
rect 11330 7060 11390 7080
rect 11440 8240 11500 8260
rect 11440 7080 11450 8240
rect 11490 7080 11500 8240
rect 11440 6990 11500 7080
rect 11550 8240 11610 8430
rect 11550 7080 11560 8240
rect 11600 7080 11610 8240
rect 11550 7060 11610 7080
rect 11660 8240 11720 8260
rect 11660 7080 11670 8240
rect 11710 7080 11720 8240
rect 11660 6990 11720 7080
rect 11770 8240 11830 8430
rect 11770 7080 11780 8240
rect 11820 7080 11830 8240
rect 11770 7060 11830 7080
rect 11880 8240 11940 8260
rect 11880 7080 11890 8240
rect 11930 7080 11940 8240
rect 11880 6990 11940 7080
rect 11990 8240 12050 8430
rect 11990 7080 12000 8240
rect 12040 7080 12050 8240
rect 11990 7060 12050 7080
rect 12100 8240 12160 8260
rect 12100 7080 12110 8240
rect 12150 7080 12160 8240
rect 12100 6990 12160 7080
rect 12210 8240 12270 8430
rect 12210 7080 12220 8240
rect 12260 7080 12270 8240
rect 12210 7060 12270 7080
rect 12320 8240 12380 8260
rect 12320 7080 12330 8240
rect 12370 7080 12380 8240
rect 12320 6990 12380 7080
rect 12430 8240 12490 8430
rect 12430 7080 12440 8240
rect 12480 7080 12490 8240
rect 12430 7060 12490 7080
rect 12540 8240 12600 8260
rect 12540 7080 12550 8240
rect 12590 7080 12600 8240
rect 12540 6990 12600 7080
rect 12650 8240 12710 8430
rect 12650 7080 12660 8240
rect 12700 7080 12710 8240
rect 12650 7060 12710 7080
rect 12760 8240 12820 8260
rect 12760 7080 12770 8240
rect 12810 7080 12820 8240
rect 12760 6990 12820 7080
rect 12870 8240 12930 8430
rect 12870 7080 12880 8240
rect 12920 7080 12930 8240
rect 12870 7060 12930 7080
rect 12980 8240 13040 8260
rect 12980 7080 12990 8240
rect 13030 7080 13040 8240
rect 12980 6990 13040 7080
rect 13090 8240 13150 8430
rect 13390 8420 13430 8430
rect 13560 8480 13600 8490
rect 13560 8430 16920 8480
rect 13560 8420 13600 8430
rect 13390 8400 13600 8420
rect 13090 7080 13100 8240
rect 13140 7080 13150 8240
rect 13090 7060 13150 7080
rect 13200 8240 13260 8260
rect 13200 7080 13210 8240
rect 13250 7080 13260 8240
rect 13200 6990 13260 7080
rect 13670 8240 13730 8260
rect 13670 7080 13680 8240
rect 13720 7080 13730 8240
rect 13670 6990 13730 7080
rect 13780 8240 13840 8430
rect 13780 7080 13790 8240
rect 13830 7080 13840 8240
rect 13780 7060 13840 7080
rect 13890 8240 13950 8260
rect 13890 7080 13900 8240
rect 13940 7080 13950 8240
rect 13890 6990 13950 7080
rect 14000 8240 14060 8430
rect 14000 7080 14010 8240
rect 14050 7080 14060 8240
rect 14000 7060 14060 7080
rect 14110 8240 14170 8260
rect 14110 7080 14120 8240
rect 14160 7080 14170 8240
rect 14110 6990 14170 7080
rect 14220 8240 14280 8430
rect 14220 7080 14230 8240
rect 14270 7080 14280 8240
rect 14220 7060 14280 7080
rect 14330 8240 14390 8260
rect 14330 7080 14340 8240
rect 14380 7080 14390 8240
rect 14330 6990 14390 7080
rect 14440 8240 14500 8430
rect 14440 7080 14450 8240
rect 14490 7080 14500 8240
rect 14440 7060 14500 7080
rect 14550 8240 14610 8260
rect 14550 7080 14560 8240
rect 14600 7080 14610 8240
rect 14550 6990 14610 7080
rect 14660 8240 14720 8430
rect 14660 7080 14670 8240
rect 14710 7080 14720 8240
rect 14660 7060 14720 7080
rect 14770 8240 14830 8260
rect 14770 7080 14780 8240
rect 14820 7080 14830 8240
rect 14770 6990 14830 7080
rect 14880 8240 14940 8430
rect 14880 7080 14890 8240
rect 14930 7080 14940 8240
rect 14880 7060 14940 7080
rect 14990 8240 15050 8260
rect 14990 7080 15000 8240
rect 15040 7080 15050 8240
rect 14990 6990 15050 7080
rect 15100 8240 15160 8430
rect 15100 7080 15110 8240
rect 15150 7080 15160 8240
rect 15100 7060 15160 7080
rect 15210 8240 15270 8260
rect 15210 7080 15220 8240
rect 15260 7080 15270 8240
rect 15210 6990 15270 7080
rect 15320 8240 15380 8430
rect 15320 7080 15330 8240
rect 15370 7080 15380 8240
rect 15320 7060 15380 7080
rect 15430 8240 15490 8260
rect 15430 7080 15440 8240
rect 15480 7080 15490 8240
rect 15430 6990 15490 7080
rect 15540 8240 15600 8430
rect 15540 7080 15550 8240
rect 15590 7080 15600 8240
rect 15540 7060 15600 7080
rect 15650 8240 15710 8260
rect 15650 7080 15660 8240
rect 15700 7080 15710 8240
rect 15650 6990 15710 7080
rect 15760 8240 15820 8430
rect 15760 7080 15770 8240
rect 15810 7080 15820 8240
rect 15760 7060 15820 7080
rect 15870 8240 15930 8260
rect 15870 7080 15880 8240
rect 15920 7080 15930 8240
rect 15870 6990 15930 7080
rect 15980 8240 16040 8430
rect 15980 7080 15990 8240
rect 16030 7080 16040 8240
rect 15980 7060 16040 7080
rect 16090 8240 16150 8260
rect 16090 7080 16100 8240
rect 16140 7080 16150 8240
rect 16090 6990 16150 7080
rect 16200 8240 16260 8430
rect 16200 7080 16210 8240
rect 16250 7080 16260 8240
rect 16200 7060 16260 7080
rect 16310 8240 16370 8260
rect 16310 7080 16320 8240
rect 16360 7080 16370 8240
rect 16310 6990 16370 7080
rect 16420 8240 16480 8430
rect 16420 7080 16430 8240
rect 16470 7080 16480 8240
rect 16420 7060 16480 7080
rect 16530 8240 16590 8260
rect 16530 7080 16540 8240
rect 16580 7080 16590 8240
rect 16530 6990 16590 7080
rect 16640 8240 16700 8430
rect 16640 7080 16650 8240
rect 16690 7080 16700 8240
rect 16640 7060 16700 7080
rect 16750 8240 16810 8260
rect 16750 7080 16760 8240
rect 16800 7080 16810 8240
rect 16750 6990 16810 7080
rect 16860 8240 16920 8430
rect 17020 8360 17130 8370
rect 17020 8310 17050 8360
rect 17100 8310 17130 8360
rect 17020 8300 17130 8310
rect 16860 7080 16870 8240
rect 16910 7080 16920 8240
rect 16860 7060 16920 7080
rect 16970 8240 17030 8260
rect 16970 7080 16980 8240
rect 17020 7080 17030 8240
rect 16970 6990 17030 7080
rect 9870 6980 17060 6990
rect 9870 6930 9900 6980
rect 9960 6930 10120 6980
rect 10180 6930 10340 6980
rect 10400 6930 10560 6980
rect 10620 6930 10780 6980
rect 10840 6930 11000 6980
rect 11060 6930 11220 6980
rect 11280 6930 11440 6980
rect 11500 6930 11660 6980
rect 11720 6930 11880 6980
rect 11940 6930 12100 6980
rect 12160 6930 12320 6980
rect 12380 6930 12540 6980
rect 12600 6930 12760 6980
rect 12820 6930 12980 6980
rect 13040 6930 13200 6980
rect 13260 6930 13670 6980
rect 13730 6930 13890 6980
rect 13950 6930 14110 6980
rect 14170 6930 14330 6980
rect 14390 6930 14550 6980
rect 14610 6930 14770 6980
rect 14830 6930 14990 6980
rect 15050 6930 15210 6980
rect 15270 6930 15430 6980
rect 15490 6930 15650 6980
rect 15710 6930 15870 6980
rect 15930 6930 16090 6980
rect 16150 6930 16310 6980
rect 16370 6930 16530 6980
rect 16590 6930 16750 6980
rect 16810 6930 16970 6980
rect 17030 6930 17060 6980
rect 9870 6920 17060 6930
rect 13600 5990 17020 6000
rect 13600 5940 13630 5990
rect 13690 5940 13850 5990
rect 13910 5940 14070 5990
rect 14130 5940 14290 5990
rect 14350 5940 14510 5990
rect 14570 5940 14730 5990
rect 14790 5940 14950 5990
rect 15010 5940 15170 5990
rect 15230 5940 15390 5990
rect 15450 5940 15610 5990
rect 15670 5940 15830 5990
rect 15890 5940 16050 5990
rect 16110 5940 16270 5990
rect 16330 5940 16490 5990
rect 16550 5940 16710 5990
rect 16770 5940 16930 5990
rect 16990 5940 17020 5990
rect 13600 5930 17020 5940
rect 13340 5880 13550 5900
rect 9870 5870 13380 5880
rect 9870 5830 9930 5870
rect 9970 5830 10010 5870
rect 10050 5830 10090 5870
rect 10130 5830 10170 5870
rect 10210 5830 10250 5870
rect 10290 5830 10330 5870
rect 10370 5830 10410 5870
rect 10450 5830 10490 5870
rect 10530 5830 10610 5870
rect 10650 5830 10690 5870
rect 10730 5830 10770 5870
rect 10810 5830 10850 5870
rect 10890 5830 10930 5870
rect 10970 5830 11010 5870
rect 11050 5830 11090 5870
rect 11130 5830 11170 5870
rect 11210 5830 11250 5870
rect 11290 5830 11370 5870
rect 11410 5830 11450 5870
rect 11490 5830 11530 5870
rect 11570 5830 11610 5870
rect 11650 5830 11690 5870
rect 11730 5830 11770 5870
rect 11810 5830 11850 5870
rect 11890 5830 11930 5870
rect 11970 5830 12010 5870
rect 12050 5830 12130 5870
rect 12170 5830 12210 5870
rect 12250 5830 12290 5870
rect 12330 5830 12370 5870
rect 12410 5830 12450 5870
rect 12490 5830 12530 5870
rect 12570 5830 12610 5870
rect 12650 5830 12690 5870
rect 12730 5830 12770 5870
rect 12810 5830 12850 5870
rect 12890 5830 12930 5870
rect 12970 5830 13010 5870
rect 13050 5830 13090 5870
rect 13130 5830 13380 5870
rect 9870 5820 13380 5830
rect 13510 5820 13550 5880
rect 9870 5600 9930 5820
rect 9870 4440 9880 5600
rect 9920 4440 9930 5600
rect 9870 4420 9930 4440
rect 9980 5600 10040 5620
rect 9980 4440 9990 5600
rect 10030 4440 10040 5600
rect 9840 4140 9940 4160
rect 9840 4070 9850 4140
rect 9930 4130 9940 4140
rect 9980 4130 10040 4440
rect 10090 5600 10150 5820
rect 10090 4440 10100 5600
rect 10140 4440 10150 5600
rect 10090 4420 10150 4440
rect 10200 5600 10260 5620
rect 10200 4440 10210 5600
rect 10250 4440 10260 5600
rect 10200 4130 10260 4440
rect 10310 5600 10370 5820
rect 10310 4440 10320 5600
rect 10360 4440 10370 5600
rect 10310 4420 10370 4440
rect 10420 5600 10480 5620
rect 10420 4440 10430 5600
rect 10470 4440 10480 5600
rect 10420 4130 10480 4440
rect 10530 5600 10590 5820
rect 10530 4440 10540 5600
rect 10580 4440 10590 5600
rect 10530 4420 10590 4440
rect 10640 5600 10700 5620
rect 10640 4440 10650 5600
rect 10690 4440 10700 5600
rect 10640 4130 10700 4440
rect 10750 5600 10810 5820
rect 10750 4440 10760 5600
rect 10800 4440 10810 5600
rect 10750 4420 10810 4440
rect 10860 5600 10920 5620
rect 10860 4440 10870 5600
rect 10910 4440 10920 5600
rect 10860 4130 10920 4440
rect 10970 5600 11030 5820
rect 10970 4440 10980 5600
rect 11020 4440 11030 5600
rect 10970 4420 11030 4440
rect 11080 5600 11140 5620
rect 11080 4440 11090 5600
rect 11130 4440 11140 5600
rect 11080 4130 11140 4440
rect 11190 5600 11250 5820
rect 11190 4440 11200 5600
rect 11240 4440 11250 5600
rect 11190 4420 11250 4440
rect 11300 5600 11360 5620
rect 11300 4440 11310 5600
rect 11350 4440 11360 5600
rect 11300 4130 11360 4440
rect 11410 5600 11470 5820
rect 11410 4440 11420 5600
rect 11460 4440 11470 5600
rect 11410 4420 11470 4440
rect 11520 5600 11580 5620
rect 11520 4440 11530 5600
rect 11570 4440 11580 5600
rect 11520 4130 11580 4440
rect 11630 5600 11690 5820
rect 11630 4440 11640 5600
rect 11680 4440 11690 5600
rect 11630 4420 11690 4440
rect 11740 5600 11800 5620
rect 11740 4440 11750 5600
rect 11790 4440 11800 5600
rect 11740 4130 11800 4440
rect 11850 5600 11910 5820
rect 11850 4440 11860 5600
rect 11900 4440 11910 5600
rect 11850 4420 11910 4440
rect 11960 5600 12020 5620
rect 11960 4440 11970 5600
rect 12010 4440 12020 5600
rect 11960 4130 12020 4440
rect 12070 5600 12130 5820
rect 12070 4440 12080 5600
rect 12120 4440 12130 5600
rect 12070 4420 12130 4440
rect 12180 5600 12240 5620
rect 12180 4440 12190 5600
rect 12230 4440 12240 5600
rect 12180 4130 12240 4440
rect 12290 5600 12350 5820
rect 12290 4440 12300 5600
rect 12340 4440 12350 5600
rect 12290 4420 12350 4440
rect 12400 5600 12460 5620
rect 12400 4440 12410 5600
rect 12450 4440 12460 5600
rect 12400 4130 12460 4440
rect 12510 5600 12570 5820
rect 12510 4440 12520 5600
rect 12560 4440 12570 5600
rect 12510 4420 12570 4440
rect 12620 5600 12680 5620
rect 12620 4440 12630 5600
rect 12670 4440 12680 5600
rect 12620 4130 12680 4440
rect 12730 5600 12790 5820
rect 12730 4440 12740 5600
rect 12780 4440 12790 5600
rect 12730 4420 12790 4440
rect 12840 5600 12900 5620
rect 12840 4440 12850 5600
rect 12890 4440 12900 5600
rect 12840 4130 12900 4440
rect 12950 5600 13010 5820
rect 12950 4440 12960 5600
rect 13000 4440 13010 5600
rect 12950 4420 13010 4440
rect 13060 5600 13120 5620
rect 13060 4440 13070 5600
rect 13110 4440 13120 5600
rect 13060 4130 13120 4440
rect 13170 5600 13230 5820
rect 13340 5800 13550 5820
rect 13630 5840 13690 5930
rect 13170 4440 13180 5600
rect 13220 4440 13230 5600
rect 13630 4680 13640 5840
rect 13680 4680 13690 5840
rect 13630 4660 13690 4680
rect 13740 5840 13800 5860
rect 13740 4680 13750 5840
rect 13790 4680 13800 5840
rect 13170 4420 13230 4440
rect 13340 4500 13550 4520
rect 13340 4440 13380 4500
rect 13510 4490 13550 4500
rect 13740 4490 13800 4680
rect 13850 5840 13910 5930
rect 13850 4680 13860 5840
rect 13900 4680 13910 5840
rect 13850 4660 13910 4680
rect 13960 5840 14020 5860
rect 13960 4680 13970 5840
rect 14010 4680 14020 5840
rect 13960 4490 14020 4680
rect 14070 5840 14130 5930
rect 14070 4680 14080 5840
rect 14120 4680 14130 5840
rect 14070 4660 14130 4680
rect 14180 5840 14240 5860
rect 14180 4680 14190 5840
rect 14230 4680 14240 5840
rect 14180 4490 14240 4680
rect 14290 5840 14350 5930
rect 14290 4680 14300 5840
rect 14340 4680 14350 5840
rect 14290 4660 14350 4680
rect 14400 5840 14460 5860
rect 14400 4680 14410 5840
rect 14450 4680 14460 5840
rect 14400 4490 14460 4680
rect 14510 5840 14570 5930
rect 14510 4680 14520 5840
rect 14560 4680 14570 5840
rect 14510 4660 14570 4680
rect 14620 5840 14680 5860
rect 14620 4680 14630 5840
rect 14670 4680 14680 5840
rect 14620 4490 14680 4680
rect 14730 5840 14790 5930
rect 14730 4680 14740 5840
rect 14780 4680 14790 5840
rect 14730 4660 14790 4680
rect 14840 5840 14900 5860
rect 14840 4680 14850 5840
rect 14890 4680 14900 5840
rect 14840 4490 14900 4680
rect 14950 5840 15010 5930
rect 14950 4680 14960 5840
rect 15000 4680 15010 5840
rect 14950 4660 15010 4680
rect 15060 5840 15120 5860
rect 15060 4680 15070 5840
rect 15110 4680 15120 5840
rect 15060 4490 15120 4680
rect 15170 5840 15230 5930
rect 15170 4680 15180 5840
rect 15220 4680 15230 5840
rect 15170 4660 15230 4680
rect 15280 5840 15340 5860
rect 15280 4680 15290 5840
rect 15330 4680 15340 5840
rect 15280 4490 15340 4680
rect 15390 5840 15450 5930
rect 15390 4680 15400 5840
rect 15440 4680 15450 5840
rect 15390 4660 15450 4680
rect 15500 5840 15560 5860
rect 15500 4680 15510 5840
rect 15550 4680 15560 5840
rect 15500 4490 15560 4680
rect 15610 5840 15670 5930
rect 15610 4680 15620 5840
rect 15660 4680 15670 5840
rect 15610 4660 15670 4680
rect 15720 5840 15780 5860
rect 15720 4680 15730 5840
rect 15770 4680 15780 5840
rect 15720 4490 15780 4680
rect 15830 5840 15890 5930
rect 15830 4680 15840 5840
rect 15880 4680 15890 5840
rect 15830 4660 15890 4680
rect 15940 5840 16000 5860
rect 15940 4680 15950 5840
rect 15990 4680 16000 5840
rect 15940 4490 16000 4680
rect 16050 5840 16110 5930
rect 16050 4680 16060 5840
rect 16100 4680 16110 5840
rect 16050 4660 16110 4680
rect 16160 5840 16220 5860
rect 16160 4680 16170 5840
rect 16210 4680 16220 5840
rect 16160 4490 16220 4680
rect 16270 5840 16330 5930
rect 16270 4680 16280 5840
rect 16320 4680 16330 5840
rect 16270 4660 16330 4680
rect 16380 5840 16440 5860
rect 16380 4680 16390 5840
rect 16430 4680 16440 5840
rect 16380 4490 16440 4680
rect 16490 5840 16550 5930
rect 16490 4680 16500 5840
rect 16540 4680 16550 5840
rect 16490 4660 16550 4680
rect 16600 5840 16660 5860
rect 16600 4680 16610 5840
rect 16650 4680 16660 5840
rect 16600 4490 16660 4680
rect 16710 5840 16770 5930
rect 16710 4680 16720 5840
rect 16760 4680 16770 5840
rect 16710 4660 16770 4680
rect 16820 5840 16880 5860
rect 16820 4680 16830 5840
rect 16870 4680 16880 5840
rect 16820 4490 16880 4680
rect 16930 5840 16990 5930
rect 16930 4680 16940 5840
rect 16980 4680 16990 5840
rect 16930 4660 16990 4680
rect 13510 4440 16880 4490
rect 16920 4470 17030 4480
rect 13340 4420 13550 4440
rect 16920 4420 16950 4470
rect 17000 4420 17030 4470
rect 16920 4410 17030 4420
rect 13340 4340 13550 4360
rect 13340 4280 13380 4340
rect 13510 4330 13550 4340
rect 13510 4280 16880 4330
rect 13340 4260 13550 4280
rect 9930 4080 13120 4130
rect 9930 4070 9940 4080
rect 9840 4050 9940 4070
rect 9870 3790 9930 3810
rect 9870 3230 9880 3790
rect 9920 3230 9930 3790
rect 9870 3080 9930 3230
rect 9980 3790 10040 4080
rect 9980 3230 9990 3790
rect 10030 3230 10040 3790
rect 9980 3210 10040 3230
rect 10090 3790 10150 3810
rect 10090 3230 10100 3790
rect 10140 3230 10150 3790
rect 10090 3080 10150 3230
rect 10200 3790 10260 4080
rect 10200 3230 10210 3790
rect 10250 3230 10260 3790
rect 10200 3210 10260 3230
rect 10310 3790 10370 3810
rect 10310 3230 10320 3790
rect 10360 3230 10370 3790
rect 10310 3080 10370 3230
rect 10420 3790 10480 4080
rect 10420 3230 10430 3790
rect 10470 3230 10480 3790
rect 10420 3210 10480 3230
rect 10530 3790 10590 3810
rect 10530 3230 10540 3790
rect 10580 3230 10590 3790
rect 10530 3080 10590 3230
rect 10640 3790 10700 4080
rect 10640 3230 10650 3790
rect 10690 3230 10700 3790
rect 10640 3210 10700 3230
rect 10750 3790 10810 3810
rect 10750 3230 10760 3790
rect 10800 3230 10810 3790
rect 10750 3080 10810 3230
rect 10860 3790 10920 4080
rect 10860 3230 10870 3790
rect 10910 3230 10920 3790
rect 10860 3210 10920 3230
rect 10970 3790 11030 3810
rect 10970 3230 10980 3790
rect 11020 3230 11030 3790
rect 10970 3080 11030 3230
rect 11080 3790 11140 4080
rect 11080 3230 11090 3790
rect 11130 3230 11140 3790
rect 11080 3210 11140 3230
rect 11190 3790 11250 3810
rect 11190 3230 11200 3790
rect 11240 3230 11250 3790
rect 11190 3080 11250 3230
rect 11300 3790 11360 4080
rect 11300 3230 11310 3790
rect 11350 3230 11360 3790
rect 11300 3210 11360 3230
rect 11410 3790 11470 3810
rect 11410 3230 11420 3790
rect 11460 3230 11470 3790
rect 11410 3080 11470 3230
rect 11520 3790 11580 4080
rect 11520 3230 11530 3790
rect 11570 3230 11580 3790
rect 11520 3210 11580 3230
rect 11630 3790 11690 3810
rect 11630 3230 11640 3790
rect 11680 3230 11690 3790
rect 11630 3080 11690 3230
rect 11740 3790 11800 4080
rect 11740 3230 11750 3790
rect 11790 3230 11800 3790
rect 11740 3210 11800 3230
rect 11850 3790 11910 3810
rect 11850 3230 11860 3790
rect 11900 3230 11910 3790
rect 11850 3080 11910 3230
rect 11960 3790 12020 4080
rect 11960 3230 11970 3790
rect 12010 3230 12020 3790
rect 11960 3210 12020 3230
rect 12070 3790 12130 3810
rect 12070 3230 12080 3790
rect 12120 3230 12130 3790
rect 12070 3080 12130 3230
rect 12180 3790 12240 4080
rect 12180 3230 12190 3790
rect 12230 3230 12240 3790
rect 12180 3210 12240 3230
rect 12290 3790 12350 3810
rect 12290 3230 12300 3790
rect 12340 3230 12350 3790
rect 12290 3080 12350 3230
rect 12400 3790 12460 4080
rect 12400 3230 12410 3790
rect 12450 3230 12460 3790
rect 12400 3210 12460 3230
rect 12510 3790 12570 3810
rect 12510 3230 12520 3790
rect 12560 3230 12570 3790
rect 12510 3080 12570 3230
rect 12620 3790 12680 4080
rect 12620 3230 12630 3790
rect 12670 3230 12680 3790
rect 12620 3210 12680 3230
rect 12730 3790 12790 3810
rect 12730 3230 12740 3790
rect 12780 3230 12790 3790
rect 12730 3080 12790 3230
rect 12840 3790 12900 4080
rect 12840 3230 12850 3790
rect 12890 3230 12900 3790
rect 12840 3210 12900 3230
rect 12950 3790 13010 3810
rect 12950 3230 12960 3790
rect 13000 3230 13010 3790
rect 12950 3080 13010 3230
rect 13060 3790 13120 4080
rect 13160 4150 13270 4170
rect 13160 4090 13180 4150
rect 13250 4090 13270 4150
rect 13160 4070 13270 4090
rect 13630 4120 13690 4140
rect 13160 3960 13270 3980
rect 13160 3900 13180 3960
rect 13250 3900 13270 3960
rect 13160 3880 13270 3900
rect 13060 3230 13070 3790
rect 13110 3230 13120 3790
rect 13060 3210 13120 3230
rect 13170 3790 13230 3810
rect 13170 3230 13180 3790
rect 13220 3230 13230 3790
rect 13170 3080 13230 3230
rect 13630 3560 13640 4120
rect 13680 3560 13690 4120
rect 13630 3370 13690 3560
rect 13740 4120 13800 4280
rect 13740 3560 13750 4120
rect 13790 3560 13800 4120
rect 13740 3540 13800 3560
rect 13850 4120 13910 4140
rect 13850 3560 13860 4120
rect 13900 3560 13910 4120
rect 13850 3370 13910 3560
rect 13960 4120 14020 4280
rect 13960 3560 13970 4120
rect 14010 3560 14020 4120
rect 13960 3540 14020 3560
rect 14070 4120 14130 4140
rect 14070 3560 14080 4120
rect 14120 3560 14130 4120
rect 14070 3370 14130 3560
rect 14180 4120 14240 4280
rect 14180 3560 14190 4120
rect 14230 3560 14240 4120
rect 14180 3540 14240 3560
rect 14290 4120 14350 4140
rect 14290 3560 14300 4120
rect 14340 3560 14350 4120
rect 14290 3370 14350 3560
rect 14400 4120 14460 4280
rect 14400 3560 14410 4120
rect 14450 3560 14460 4120
rect 14400 3540 14460 3560
rect 14510 4120 14570 4140
rect 14510 3560 14520 4120
rect 14560 3560 14570 4120
rect 14510 3370 14570 3560
rect 14620 4120 14680 4280
rect 14620 3560 14630 4120
rect 14670 3560 14680 4120
rect 14620 3540 14680 3560
rect 14730 4120 14790 4140
rect 14730 3560 14740 4120
rect 14780 3560 14790 4120
rect 14730 3370 14790 3560
rect 14840 4120 14900 4280
rect 14840 3560 14850 4120
rect 14890 3560 14900 4120
rect 14840 3540 14900 3560
rect 14950 4120 15010 4140
rect 14950 3560 14960 4120
rect 15000 3560 15010 4120
rect 14950 3370 15010 3560
rect 15060 4120 15120 4280
rect 15060 3560 15070 4120
rect 15110 3560 15120 4120
rect 15060 3540 15120 3560
rect 15170 4120 15230 4140
rect 15170 3560 15180 4120
rect 15220 3560 15230 4120
rect 15170 3370 15230 3560
rect 15280 4120 15340 4280
rect 15280 3560 15290 4120
rect 15330 3560 15340 4120
rect 15280 3540 15340 3560
rect 15390 4120 15450 4140
rect 15390 3560 15400 4120
rect 15440 3560 15450 4120
rect 15390 3370 15450 3560
rect 15500 4120 15560 4280
rect 15500 3560 15510 4120
rect 15550 3560 15560 4120
rect 15500 3540 15560 3560
rect 15610 4120 15670 4140
rect 15610 3560 15620 4120
rect 15660 3560 15670 4120
rect 15610 3370 15670 3560
rect 15720 4120 15780 4280
rect 15720 3560 15730 4120
rect 15770 3560 15780 4120
rect 15720 3540 15780 3560
rect 15830 4120 15890 4140
rect 15830 3560 15840 4120
rect 15880 3560 15890 4120
rect 15830 3370 15890 3560
rect 15940 4120 16000 4280
rect 15940 3560 15950 4120
rect 15990 3560 16000 4120
rect 15940 3540 16000 3560
rect 16050 4120 16110 4140
rect 16050 3560 16060 4120
rect 16100 3560 16110 4120
rect 16050 3370 16110 3560
rect 16160 4120 16220 4280
rect 16160 3560 16170 4120
rect 16210 3560 16220 4120
rect 16160 3540 16220 3560
rect 16270 4120 16330 4140
rect 16270 3560 16280 4120
rect 16320 3560 16330 4120
rect 16270 3370 16330 3560
rect 16380 4120 16440 4280
rect 16380 3560 16390 4120
rect 16430 3560 16440 4120
rect 16380 3540 16440 3560
rect 16490 4120 16550 4140
rect 16490 3560 16500 4120
rect 16540 3560 16550 4120
rect 16490 3370 16550 3560
rect 16600 4120 16660 4280
rect 16600 3560 16610 4120
rect 16650 3560 16660 4120
rect 16600 3540 16660 3560
rect 16710 4120 16770 4140
rect 16710 3560 16720 4120
rect 16760 3560 16770 4120
rect 16710 3370 16770 3560
rect 16820 4120 16880 4280
rect 16820 3560 16830 4120
rect 16870 3560 16880 4120
rect 16820 3540 16880 3560
rect 16930 4120 16990 4140
rect 16930 3560 16940 4120
rect 16980 3560 16990 4120
rect 16930 3370 16990 3560
rect 13630 3320 16990 3370
rect 13280 3080 13490 3100
rect 9870 3020 13320 3080
rect 13450 3020 13490 3080
rect 13280 3000 13490 3020
rect 13630 3010 13690 3320
rect 13850 3010 13910 3320
rect 14070 3010 14130 3320
rect 14290 3010 14350 3320
rect 14510 3010 14570 3320
rect 14730 3010 14790 3320
rect 14950 3010 15010 3320
rect 15170 3010 15230 3320
rect 15390 3010 15450 3320
rect 15610 3010 15670 3320
rect 15830 3010 15890 3320
rect 16050 3010 16110 3320
rect 16270 3010 16330 3320
rect 16490 3010 16550 3320
rect 16710 3010 16770 3320
rect 16920 3240 17020 3250
rect 16920 3190 16950 3240
rect 17000 3190 17020 3240
rect 16920 3180 17020 3190
rect 13600 3000 17020 3010
rect 13600 2950 13630 3000
rect 13690 2950 13850 3000
rect 13910 2950 14070 3000
rect 14130 2950 14290 3000
rect 14350 2950 14510 3000
rect 14570 2950 14730 3000
rect 14790 2950 14950 3000
rect 15010 2950 15170 3000
rect 15230 2950 15390 3000
rect 15450 2950 15610 3000
rect 15670 2950 15830 3000
rect 15890 2950 16050 3000
rect 16110 2950 16270 3000
rect 16330 2950 16490 3000
rect 16550 2950 16710 3000
rect 16770 2950 17020 3000
rect 13600 2940 17020 2950
rect 24210 2720 24290 2770
rect 24210 2660 24220 2720
rect 24280 2660 24290 2720
rect 24350 2760 25550 2770
rect 24350 2720 24370 2760
rect 25330 2720 25550 2760
rect 24350 2710 25550 2720
rect 24210 2650 25350 2660
rect 24210 2620 24370 2650
rect 24210 2560 24220 2620
rect 24280 2610 24370 2620
rect 25330 2610 25350 2650
rect 24280 2600 25350 2610
rect 24280 2560 24290 2600
rect 24210 2520 24290 2560
rect 25470 2550 25550 2710
rect 25710 2760 25780 2780
rect 25710 2720 25720 2760
rect 25770 2720 25780 2760
rect 25710 2700 25780 2720
rect 25710 2640 25780 2660
rect 25710 2600 25720 2640
rect 25770 2600 25780 2640
rect 25710 2580 25780 2600
rect 24210 2460 24220 2520
rect 24280 2460 24290 2520
rect 24350 2540 25550 2550
rect 24350 2500 24370 2540
rect 25330 2500 25550 2540
rect 24350 2490 25550 2500
rect 24210 2440 24290 2460
rect 24210 2430 25350 2440
rect 24210 2420 24370 2430
rect 24210 2360 24220 2420
rect 24280 2390 24370 2420
rect 25330 2390 25350 2430
rect 24280 2380 25350 2390
rect 24280 2360 24290 2380
rect 24210 2320 24290 2360
rect 25470 2330 25550 2490
rect 25710 2520 25780 2540
rect 25710 2480 25720 2520
rect 25770 2480 25780 2520
rect 25710 2460 25780 2480
rect 25710 2400 25780 2420
rect 25710 2360 25720 2400
rect 25770 2360 25780 2400
rect 25710 2340 25780 2360
rect 24210 2260 24220 2320
rect 24280 2260 24290 2320
rect 24350 2320 25550 2330
rect 24350 2280 24370 2320
rect 25330 2280 25550 2320
rect 24350 2270 25550 2280
rect 24210 2220 24290 2260
rect 24210 2160 24220 2220
rect 24280 2210 25350 2220
rect 24280 2170 24370 2210
rect 25330 2170 25350 2210
rect 24280 2160 25350 2170
rect 24210 2120 24290 2160
rect 24210 2060 24220 2120
rect 24280 2060 24290 2120
rect 25470 2110 25550 2270
rect 25710 2280 25780 2300
rect 25710 2240 25720 2280
rect 25770 2240 25780 2280
rect 25710 2220 25780 2240
rect 24210 2030 24290 2060
rect 24350 2100 25550 2110
rect 25710 2160 25780 2180
rect 25710 2120 25720 2160
rect 25770 2120 25780 2160
rect 25710 2100 25780 2120
rect 24350 2060 24370 2100
rect 25330 2060 25550 2100
rect 24350 2050 25550 2060
rect 25470 1970 25550 2050
rect 9850 1920 17020 1930
rect 9850 1870 9890 1920
rect 9950 1870 10110 1920
rect 10170 1870 10330 1920
rect 10390 1870 10550 1920
rect 10610 1870 10770 1920
rect 10830 1870 10990 1920
rect 11050 1870 11210 1920
rect 11270 1870 11430 1920
rect 11490 1870 11650 1920
rect 11710 1870 11870 1920
rect 11930 1870 12090 1920
rect 12150 1870 12310 1920
rect 12370 1870 12530 1920
rect 12590 1870 12750 1920
rect 12810 1870 12970 1920
rect 13030 1870 13630 1920
rect 13690 1870 13850 1920
rect 13910 1870 14070 1920
rect 14130 1870 14290 1920
rect 14350 1870 14510 1920
rect 14570 1870 14730 1920
rect 14790 1870 14950 1920
rect 15010 1870 15170 1920
rect 15230 1870 15390 1920
rect 15450 1870 15610 1920
rect 15670 1870 15830 1920
rect 15890 1870 16050 1920
rect 16110 1870 16270 1920
rect 16330 1870 16490 1920
rect 16550 1870 16710 1920
rect 16770 1870 17020 1920
rect 9850 1860 17020 1870
rect 25470 1910 25480 1970
rect 25540 1910 25550 1970
rect 25470 1860 25550 1910
rect 9890 1550 9950 1860
rect 10110 1550 10170 1860
rect 10330 1550 10390 1860
rect 10550 1550 10610 1860
rect 10770 1550 10830 1860
rect 10990 1550 11050 1860
rect 11210 1550 11270 1860
rect 11430 1550 11490 1860
rect 11650 1550 11710 1860
rect 11870 1550 11930 1860
rect 12090 1550 12150 1860
rect 12310 1550 12370 1860
rect 12530 1550 12590 1860
rect 12750 1550 12810 1860
rect 12970 1550 13030 1860
rect 13180 1680 13280 1690
rect 13180 1630 13210 1680
rect 13260 1630 13280 1680
rect 13180 1620 13280 1630
rect 9890 1500 13250 1550
rect 9890 1310 9950 1500
rect 9890 750 9900 1310
rect 9940 750 9950 1310
rect 9890 730 9950 750
rect 10000 1310 10060 1330
rect 10000 750 10010 1310
rect 10050 750 10060 1310
rect 10000 580 10060 750
rect 10110 1310 10170 1500
rect 10110 750 10120 1310
rect 10160 750 10170 1310
rect 10110 730 10170 750
rect 10220 1310 10280 1330
rect 10220 750 10230 1310
rect 10270 750 10280 1310
rect 10220 580 10280 750
rect 10330 1310 10390 1500
rect 10330 750 10340 1310
rect 10380 750 10390 1310
rect 10330 730 10390 750
rect 10440 1310 10500 1330
rect 10440 750 10450 1310
rect 10490 750 10500 1310
rect 10440 580 10500 750
rect 10550 1310 10610 1500
rect 10550 750 10560 1310
rect 10600 750 10610 1310
rect 10550 730 10610 750
rect 10660 1310 10720 1330
rect 10660 750 10670 1310
rect 10710 750 10720 1310
rect 10660 580 10720 750
rect 10770 1310 10830 1500
rect 10770 750 10780 1310
rect 10820 750 10830 1310
rect 10770 730 10830 750
rect 10880 1310 10940 1330
rect 10880 750 10890 1310
rect 10930 750 10940 1310
rect 10880 580 10940 750
rect 10990 1310 11050 1500
rect 10990 750 11000 1310
rect 11040 750 11050 1310
rect 10990 730 11050 750
rect 11100 1310 11160 1330
rect 11100 750 11110 1310
rect 11150 750 11160 1310
rect 11100 580 11160 750
rect 11210 1310 11270 1500
rect 11210 750 11220 1310
rect 11260 750 11270 1310
rect 11210 730 11270 750
rect 11320 1310 11380 1330
rect 11320 750 11330 1310
rect 11370 750 11380 1310
rect 11320 580 11380 750
rect 11430 1310 11490 1500
rect 11430 750 11440 1310
rect 11480 750 11490 1310
rect 11430 730 11490 750
rect 11540 1310 11600 1330
rect 11540 750 11550 1310
rect 11590 750 11600 1310
rect 11540 580 11600 750
rect 11650 1310 11710 1500
rect 11650 750 11660 1310
rect 11700 750 11710 1310
rect 11650 730 11710 750
rect 11760 1310 11820 1330
rect 11760 750 11770 1310
rect 11810 750 11820 1310
rect 11760 580 11820 750
rect 11870 1310 11930 1500
rect 11870 750 11880 1310
rect 11920 750 11930 1310
rect 11870 730 11930 750
rect 11980 1310 12040 1330
rect 11980 750 11990 1310
rect 12030 750 12040 1310
rect 11980 580 12040 750
rect 12090 1310 12150 1500
rect 12090 750 12100 1310
rect 12140 750 12150 1310
rect 12090 730 12150 750
rect 12200 1310 12260 1330
rect 12200 750 12210 1310
rect 12250 750 12260 1310
rect 12200 580 12260 750
rect 12310 1310 12370 1500
rect 12310 750 12320 1310
rect 12360 750 12370 1310
rect 12310 730 12370 750
rect 12420 1310 12480 1330
rect 12420 750 12430 1310
rect 12470 750 12480 1310
rect 12420 580 12480 750
rect 12530 1310 12590 1500
rect 12530 750 12540 1310
rect 12580 750 12590 1310
rect 12530 730 12590 750
rect 12640 1310 12700 1330
rect 12640 750 12650 1310
rect 12690 750 12700 1310
rect 12640 580 12700 750
rect 12750 1310 12810 1500
rect 12750 750 12760 1310
rect 12800 750 12810 1310
rect 12750 730 12810 750
rect 12860 1310 12920 1330
rect 12860 750 12870 1310
rect 12910 750 12920 1310
rect 12860 580 12920 750
rect 12970 1310 13030 1500
rect 12970 750 12980 1310
rect 13020 750 13030 1310
rect 12970 730 13030 750
rect 13080 1310 13140 1330
rect 13080 750 13090 1310
rect 13130 750 13140 1310
rect 13080 580 13140 750
rect 13190 1310 13250 1500
rect 13190 750 13200 1310
rect 13240 750 13250 1310
rect 13190 730 13250 750
rect 13630 1540 13690 1860
rect 13850 1540 13910 1860
rect 14070 1540 14130 1860
rect 14290 1540 14350 1860
rect 14510 1540 14570 1860
rect 14730 1540 14790 1860
rect 14950 1540 15010 1860
rect 15170 1540 15230 1860
rect 15390 1540 15450 1860
rect 15610 1540 15670 1860
rect 15830 1540 15890 1860
rect 16050 1540 16110 1860
rect 16270 1540 16330 1860
rect 16490 1540 16550 1860
rect 16710 1540 16770 1860
rect 13630 1490 16990 1540
rect 13630 1300 13690 1490
rect 13630 740 13640 1300
rect 13680 740 13690 1300
rect 13630 720 13690 740
rect 13740 1300 13800 1320
rect 13740 740 13750 1300
rect 13790 740 13800 1300
rect 13320 600 13530 620
rect 13320 580 13360 600
rect 9870 530 13360 580
rect 13490 580 13530 600
rect 13740 580 13800 740
rect 13850 1300 13910 1490
rect 13850 740 13860 1300
rect 13900 740 13910 1300
rect 13850 720 13910 740
rect 13960 1300 14020 1320
rect 13960 740 13970 1300
rect 14010 740 14020 1300
rect 13960 580 14020 740
rect 14070 1300 14130 1490
rect 14070 740 14080 1300
rect 14120 740 14130 1300
rect 14070 720 14130 740
rect 14180 1300 14240 1320
rect 14180 740 14190 1300
rect 14230 740 14240 1300
rect 14180 580 14240 740
rect 14290 1300 14350 1490
rect 14290 740 14300 1300
rect 14340 740 14350 1300
rect 14290 720 14350 740
rect 14400 1300 14460 1320
rect 14400 740 14410 1300
rect 14450 740 14460 1300
rect 14400 580 14460 740
rect 14510 1300 14570 1490
rect 14510 740 14520 1300
rect 14560 740 14570 1300
rect 14510 720 14570 740
rect 14620 1300 14680 1320
rect 14620 740 14630 1300
rect 14670 740 14680 1300
rect 14620 580 14680 740
rect 14730 1300 14790 1490
rect 14730 740 14740 1300
rect 14780 740 14790 1300
rect 14730 720 14790 740
rect 14840 1300 14900 1320
rect 14840 740 14850 1300
rect 14890 740 14900 1300
rect 14840 580 14900 740
rect 14950 1300 15010 1490
rect 14950 740 14960 1300
rect 15000 740 15010 1300
rect 14950 720 15010 740
rect 15060 1300 15120 1320
rect 15060 740 15070 1300
rect 15110 740 15120 1300
rect 15060 580 15120 740
rect 15170 1300 15230 1490
rect 15170 740 15180 1300
rect 15220 740 15230 1300
rect 15170 720 15230 740
rect 15280 1300 15340 1320
rect 15280 740 15290 1300
rect 15330 740 15340 1300
rect 15280 580 15340 740
rect 15390 1300 15450 1490
rect 15390 740 15400 1300
rect 15440 740 15450 1300
rect 15390 720 15450 740
rect 15500 1300 15560 1320
rect 15500 740 15510 1300
rect 15550 740 15560 1300
rect 15500 580 15560 740
rect 15610 1300 15670 1490
rect 15610 740 15620 1300
rect 15660 740 15670 1300
rect 15610 720 15670 740
rect 15720 1300 15780 1320
rect 15720 740 15730 1300
rect 15770 740 15780 1300
rect 15720 580 15780 740
rect 15830 1300 15890 1490
rect 15830 740 15840 1300
rect 15880 740 15890 1300
rect 15830 720 15890 740
rect 15940 1300 16000 1320
rect 15940 740 15950 1300
rect 15990 740 16000 1300
rect 15940 580 16000 740
rect 16050 1300 16110 1490
rect 16050 740 16060 1300
rect 16100 740 16110 1300
rect 16050 720 16110 740
rect 16160 1300 16220 1320
rect 16160 740 16170 1300
rect 16210 740 16220 1300
rect 16160 580 16220 740
rect 16270 1300 16330 1490
rect 16270 740 16280 1300
rect 16320 740 16330 1300
rect 16270 720 16330 740
rect 16380 1300 16440 1320
rect 16380 740 16390 1300
rect 16430 740 16440 1300
rect 16380 580 16440 740
rect 16490 1300 16550 1490
rect 16490 740 16500 1300
rect 16540 740 16550 1300
rect 16490 720 16550 740
rect 16600 1300 16660 1320
rect 16600 740 16610 1300
rect 16650 740 16660 1300
rect 16600 580 16660 740
rect 16710 1300 16770 1490
rect 16710 740 16720 1300
rect 16760 740 16770 1300
rect 16710 720 16770 740
rect 16820 1300 16880 1320
rect 16820 740 16830 1300
rect 16870 740 16880 1300
rect 16820 580 16880 740
rect 16930 1300 16990 1490
rect 17030 1420 17130 1430
rect 17030 1370 17060 1420
rect 17110 1370 17130 1420
rect 17030 1360 17130 1370
rect 16930 740 16940 1300
rect 16980 740 16990 1300
rect 16930 720 16990 740
rect 13490 530 16990 580
rect 13320 510 13530 530
<< viali >>
rect 21830 43280 21890 43350
rect 21930 43280 21990 43350
rect 22030 43280 22090 43350
rect 22130 43280 22190 43350
rect 22230 43280 22290 43350
rect 22330 43280 22390 43350
rect 22430 43280 22490 43350
rect 22530 43280 22590 43350
rect 22630 43280 22690 43350
rect 22730 43280 22790 43350
rect 22830 43280 22890 43350
rect 22930 43280 22990 43350
rect 23030 43280 23090 43350
rect 23130 43280 23190 43350
rect 23230 43280 23290 43350
rect 23330 43280 23390 43350
rect 23430 43280 23490 43350
rect 23530 43280 23590 43350
rect 2469 42110 2519 42160
rect 2559 42110 2609 42160
rect 2649 42110 2699 42160
rect 2739 42110 2789 42160
rect 2829 42110 2879 42160
rect 2919 42110 2969 42160
rect 2789 42010 2829 42050
rect 2679 41580 2719 41620
rect 3429 41900 3479 41950
rect 3519 41900 3569 41950
rect 3609 41900 3659 41950
rect 3699 41900 3749 41950
rect 3789 41900 3839 41950
rect 3879 41900 3929 41950
rect 3969 41900 4019 41950
rect 4059 41900 4109 41950
rect 4149 41900 4199 41950
rect 4239 41900 4289 41950
rect 4579 41890 4639 41950
rect 6009 41910 6069 41970
rect 6119 41910 6179 41970
rect 6229 41910 6289 41970
rect 6339 41910 6399 41970
rect 6449 41910 6509 41970
rect 6559 41910 6619 41970
rect 6669 41910 6729 41970
rect 6779 41910 6839 41970
rect 6889 41910 6949 41970
rect 6999 41910 7059 41970
rect 7109 41910 7169 41970
rect 7219 41910 7279 41970
rect 7329 41910 7389 41970
rect 7439 41910 7499 41970
rect 7549 41910 7609 41970
rect 7659 41910 7719 41970
rect 7769 41910 7829 41970
rect 7879 41910 7939 41970
rect 7989 41910 8049 41970
rect 8099 41910 8159 41970
rect 8209 41910 8269 41970
rect 8319 41910 8379 41970
rect 8429 41910 8489 41970
rect 8539 41910 8599 41970
rect 8649 41910 8709 41970
rect 8759 41910 8819 41970
rect 8869 41910 8929 41970
rect 8979 41910 9039 41970
rect 9089 41910 9149 41970
rect 9199 41910 9259 41970
rect 9309 41910 9369 41970
rect 9419 41910 9479 41970
rect 9529 41910 9589 41970
rect 9639 41910 9699 41970
rect 9749 41910 9809 41970
rect 9859 41910 9919 41970
rect 21630 41920 21700 41980
rect 22340 43090 22400 43150
rect 22070 42070 22130 42130
rect 22590 42060 22630 42100
rect 23110 42100 23150 42140
rect 23000 41990 23040 42030
rect 23470 42280 23510 42320
rect 23500 42170 23540 42210
rect 21850 41930 21890 41970
rect 22590 41930 22630 41970
rect 3089 41640 3169 41680
rect 2899 41540 2939 41580
rect 2789 41470 2829 41510
rect 3179 41460 3239 41520
rect 2989 40900 3029 40940
rect 3469 40950 3509 40990
rect 2769 40620 2809 40660
rect 2879 40730 2919 40770
rect 3099 40740 3139 40780
rect 2999 40620 3039 40660
rect 2879 40490 2919 40530
rect 2759 39650 2799 39690
rect 4419 40740 4459 40780
rect 5969 41240 6009 41280
rect 6069 41240 6109 41280
rect 5359 40940 5399 40980
rect 6199 41240 6239 41280
rect 6409 41240 6449 41280
rect 6539 41240 6579 41280
rect 6969 41240 7009 41280
rect 7099 41240 7139 41280
rect 23120 41930 23160 41970
rect 22590 41760 22630 41800
rect 7969 41240 8009 41280
rect 8159 41240 8199 41280
rect 9959 41230 10009 41280
rect 22450 41270 22510 41330
rect 23000 41870 23040 41910
rect 23640 41810 23720 41870
rect 23110 41760 23150 41800
rect 23500 41720 23540 41760
rect 23810 41630 23870 41690
rect 21620 41090 21680 41160
rect 21720 41090 21780 41160
rect 21830 41090 21890 41160
rect 21930 41090 21990 41160
rect 22030 41090 22090 41160
rect 22130 41090 22190 41160
rect 22230 41090 22290 41160
rect 22330 41090 22390 41160
rect 22430 41090 22490 41160
rect 22530 41090 22590 41160
rect 22630 41090 22690 41160
rect 22730 41090 22790 41160
rect 22830 41090 22890 41160
rect 22930 41090 22990 41160
rect 23030 41090 23090 41160
rect 23130 41090 23190 41160
rect 23230 41090 23290 41160
rect 23330 41090 23390 41160
rect 23430 41090 23490 41160
rect 23530 41090 23590 41160
rect 5509 40860 5569 40920
rect 6009 40850 6070 40910
rect 5459 40740 5499 40780
rect 3320 40610 3380 40670
rect 3430 40610 3490 40670
rect 3540 40610 3600 40670
rect 3650 40610 3710 40670
rect 3760 40610 3820 40670
rect 3870 40610 3930 40670
rect 3980 40610 4040 40670
rect 4090 40610 4150 40670
rect 3339 39660 3379 39700
rect 4659 40620 5399 40660
rect 6409 40590 6469 40650
rect 6519 40590 6579 40650
rect 6629 40590 6689 40650
rect 6739 40590 6799 40650
rect 6849 40590 6909 40650
rect 6959 40590 7019 40650
rect 7069 40590 7129 40650
rect 7179 40590 7239 40650
rect 7289 40590 7349 40650
rect 7399 40590 7459 40650
rect 7509 40590 7569 40650
rect 7619 40590 7679 40650
rect 7729 40590 7789 40650
rect 7839 40590 7899 40650
rect 7949 40590 8009 40650
rect 8059 40590 8119 40650
rect 8169 40590 8229 40650
rect 8279 40590 8339 40650
rect 8389 40590 8449 40650
rect 8499 40590 8559 40650
rect 8609 40590 8669 40650
rect 8719 40590 8779 40650
rect 8829 40590 8889 40650
rect 8939 40590 8999 40650
rect 9049 40590 9109 40650
rect 9159 40590 9219 40650
rect 9269 40590 9329 40650
rect 9379 40590 9439 40650
rect 9489 40590 9549 40650
rect 9599 40590 9659 40650
rect 9709 40590 9769 40650
rect 9819 40590 9879 40650
rect 6369 39920 6409 39960
rect 9929 39910 9979 39960
rect 5359 39660 5399 39700
rect 2649 39500 2709 39560
rect 2749 39500 2809 39560
rect 2849 39500 2909 39560
rect 2949 39500 3009 39560
rect 3049 39500 3109 39560
rect 3149 39500 3209 39560
rect 3249 39500 3309 39560
rect 3349 39500 3409 39560
rect 3449 39500 3509 39560
rect 3549 39500 3609 39560
rect 3649 39500 3709 39560
rect 3749 39500 3809 39560
rect 3849 39500 3909 39560
rect 3949 39500 4009 39560
rect 4049 39500 4109 39560
rect 4149 39500 4209 39560
rect 4249 39500 4309 39560
rect 4349 39500 4409 39560
rect 4449 39500 4509 39560
rect 4549 39500 4609 39560
rect 4649 39500 4709 39560
rect 4749 39500 4809 39560
rect 4849 39500 4909 39560
rect 4949 39500 5009 39560
rect 5049 39500 5109 39560
rect 5149 39500 5209 39560
rect 5249 39500 5309 39560
rect 6349 39500 6409 39560
rect 6449 39500 6509 39560
rect 6549 39500 6609 39560
rect 6649 39500 6709 39560
rect 6749 39500 6809 39560
rect 6849 39500 6909 39560
rect 6949 39500 7009 39560
rect 7049 39500 7109 39560
rect 7149 39500 7209 39560
rect 7249 39500 7309 39560
rect 7349 39500 7409 39560
rect 7479 39500 7539 39560
rect 7579 39500 7639 39560
rect 7679 39500 7739 39560
rect 7779 39500 7839 39560
rect 7879 39500 7939 39560
rect 7979 39500 8039 39560
rect 8079 39500 8139 39560
rect 8179 39500 8239 39560
rect 8279 39500 8339 39560
rect 8379 39500 8439 39560
rect 8479 39500 8539 39560
rect 8629 39500 8689 39560
rect 8729 39500 8789 39560
rect 8829 39500 8889 39560
rect 8929 39500 8989 39560
rect 9029 39500 9089 39560
rect 9129 39500 9189 39560
rect 9229 39500 9289 39560
rect 9329 39500 9389 39560
rect 9429 39500 9489 39560
rect 9529 39500 9589 39560
rect 9629 39500 9689 39560
rect 9739 39500 9799 39560
rect 9839 39500 9899 39560
rect 25330 38430 25400 38500
rect 25840 38430 25910 38500
rect 3810 37120 3870 37180
rect 3910 37120 3970 37180
rect 4010 37120 4070 37180
rect 4110 37120 4170 37180
rect 4210 37120 4270 37180
rect 4310 37120 4370 37180
rect 4410 37120 4470 37180
rect 4510 37120 4570 37180
rect 4610 37120 4670 37180
rect 4710 37120 4770 37180
rect 4810 37120 4870 37180
rect 4910 37120 4970 37180
rect 5010 37120 5070 37180
rect 5110 37120 5170 37180
rect 5210 37120 5270 37180
rect 5310 37120 5370 37180
rect 5410 37120 5470 37180
rect 5510 37120 5570 37180
rect 5610 37120 5670 37180
rect 5710 37120 5770 37180
rect 5810 37120 5870 37180
rect 5910 37120 5970 37180
rect 6010 37120 6070 37180
rect 6110 37120 6170 37180
rect 3760 34940 3810 34990
rect 4560 34930 4620 35000
rect 5310 34820 5360 34870
rect 5420 34820 5470 34870
rect 6380 36660 6440 36720
rect 6480 36660 6540 36720
rect 6580 36660 6640 36720
rect 6680 36660 6740 36720
rect 6780 36660 6840 36720
rect 6880 36660 6940 36720
rect 6980 36660 7040 36720
rect 7080 36660 7140 36720
rect 7180 36660 7240 36720
rect 7280 36660 7340 36720
rect 7380 36660 7440 36720
rect 7480 36660 7540 36720
rect 7580 36660 7640 36720
rect 7680 36660 7740 36720
rect 7780 36660 7840 36720
rect 7880 36660 7940 36720
rect 7980 36660 8040 36720
rect 8080 36660 8140 36720
rect 8180 36660 8240 36720
rect 8280 36660 8340 36720
rect 8380 36660 8440 36720
rect 8480 36660 8540 36720
rect 8580 36660 8640 36720
rect 8680 36660 8740 36720
rect 8780 36660 8840 36720
rect 8880 36660 8940 36720
rect 8980 36660 9040 36720
rect 9080 36660 9140 36720
rect 9180 36660 9240 36720
rect 9280 36660 9340 36720
rect 9380 36660 9440 36720
rect 9480 36660 9540 36720
rect 9580 36660 9640 36720
rect 9680 36660 9740 36720
rect 9780 36660 9840 36720
rect 9880 36660 9940 36720
rect 9980 36660 10040 36720
rect 10080 36660 10140 36720
rect 10180 36660 10240 36720
rect 10280 36660 10340 36720
rect 10380 36660 10440 36720
rect 10480 36660 10540 36720
rect 10580 36660 10640 36720
rect 10680 36660 10740 36720
rect 10780 36660 10840 36720
rect 6190 34810 6240 34860
rect 6340 34810 6380 34850
rect 8680 35370 8760 35460
rect 9060 34910 9100 34950
rect 15220 36270 15280 36340
rect 15320 36270 15380 36340
rect 15420 36270 15480 36340
rect 15520 36270 15580 36340
rect 15620 36270 15680 36340
rect 15720 36270 15780 36340
rect 15820 36270 15880 36340
rect 15920 36270 15980 36340
rect 16020 36270 16080 36340
rect 16120 36270 16180 36340
rect 16220 36270 16280 36340
rect 16320 36270 16380 36340
rect 16420 36270 16480 36340
rect 16520 36270 16580 36340
rect 16620 36270 16680 36340
rect 16720 36270 16780 36340
rect 16820 36270 16880 36340
rect 16920 36270 16980 36340
rect 17020 36270 17080 36340
rect 17120 36270 17180 36340
rect 17220 36270 17280 36340
rect 17320 36270 17380 36340
rect 17420 36270 17480 36340
rect 17520 36270 17580 36340
rect 17620 36270 17680 36340
rect 17720 36270 17780 36340
rect 17820 36270 17880 36340
rect 17920 36270 17980 36340
rect 18020 36270 18080 36340
rect 18120 36270 18180 36340
rect 18220 36270 18280 36340
rect 18320 36270 18380 36340
rect 18420 36270 18480 36340
rect 18520 36270 18580 36340
rect 18620 36270 18680 36340
rect 18720 36270 18780 36340
rect 18820 36270 18880 36340
rect 18920 36270 18980 36340
rect 19020 36270 19080 36340
rect 19120 36270 19180 36340
rect 19220 36270 19280 36340
rect 19320 36270 19380 36340
rect 19420 36270 19480 36340
rect 19520 36270 19580 36340
rect 19620 36270 19680 36340
rect 19720 36270 19780 36340
rect 19820 36270 19880 36340
rect 19920 36270 19980 36340
rect 20020 36270 20080 36340
rect 20120 36270 20180 36340
rect 20220 36270 20280 36340
rect 20320 36270 20380 36340
rect 20420 36270 20480 36340
rect 20520 36270 20580 36340
rect 20620 36270 20680 36340
rect 20720 36270 20780 36340
rect 20820 36270 20880 36340
rect 20920 36270 20980 36340
rect 21020 36270 21080 36340
rect 21120 36270 21180 36340
rect 21220 36270 21280 36340
rect 21320 36270 21380 36340
rect 21420 36270 21480 36340
rect 21520 36270 21580 36340
rect 21620 36270 21680 36340
rect 21720 36270 21780 36340
rect 21820 36270 21880 36340
rect 21920 36270 21980 36340
rect 22020 36270 22080 36340
rect 22120 36270 22180 36340
rect 22220 36270 22280 36340
rect 22320 36270 22380 36340
rect 22420 36270 22480 36340
rect 22520 36270 22580 36340
rect 22620 36270 22680 36340
rect 22720 36270 22780 36340
rect 22820 36270 22880 36340
rect 22920 36270 22980 36340
rect 23020 36270 23080 36340
rect 23120 36270 23180 36340
rect 23220 36270 23280 36340
rect 23320 36270 23380 36340
rect 23420 36270 23480 36340
rect 23520 36270 23580 36340
rect 23620 36270 23680 36340
rect 23720 36270 23780 36340
rect 23820 36270 23880 36340
rect 23920 36270 23980 36340
rect 24020 36270 24080 36340
rect 24120 36270 24180 36340
rect 24220 36270 24280 36340
rect 24320 36270 24380 36340
rect 24420 36270 24480 36340
rect 24520 36270 24580 36340
rect 24620 36270 24680 36340
rect 24720 36270 24780 36340
rect 24820 36270 24880 36340
rect 15200 36050 15300 36110
rect 15460 36070 15500 36110
rect 15570 35570 15640 35630
rect 15790 35570 15900 35630
rect 15460 35480 15500 35520
rect 16450 35430 16510 35490
rect 17140 35450 17180 35490
rect 6640 34810 6680 34850
rect 6720 34810 6760 34850
rect 7220 34800 7260 34840
rect 7300 34800 7340 34840
rect 7600 34800 7640 34840
rect 7680 34800 7720 34840
rect 7980 34800 8020 34840
rect 8060 34800 8100 34840
rect 8360 34800 8400 34840
rect 8440 34800 8480 34840
rect 8690 34800 8730 34840
rect 8800 34800 8840 34840
rect 7180 34150 7220 34190
rect 9300 34800 9340 34840
rect 9380 34800 9420 34840
rect 9680 34800 9720 34840
rect 9760 34800 9800 34840
rect 10060 34800 10100 34840
rect 10140 34800 10180 34840
rect 10440 34800 10480 34840
rect 10520 34800 10560 34840
rect 10820 34800 10860 34840
rect 17580 35450 17620 35490
rect 17720 35450 17760 35490
rect 18040 35450 18080 35490
rect 17650 35320 17690 35360
rect 17240 35240 17310 35310
rect 18520 35450 18560 35490
rect 18660 35450 18700 35490
rect 18980 35450 19020 35490
rect 18590 35320 18630 35360
rect 18270 35230 18340 35300
rect 17870 35160 17910 35200
rect 17470 34860 17510 34900
rect 18410 34860 18450 34900
rect 18700 34860 18740 34900
rect 20730 36090 20790 36170
rect 20730 35830 20790 35910
rect 19770 35450 19810 35490
rect 20020 35480 20060 35520
rect 19130 34910 19170 34950
rect 19320 34910 19360 34950
rect 19520 34910 19560 34950
rect 20210 35330 20250 35370
rect 21430 35450 21470 35490
rect 22100 35450 22140 35490
rect 18310 34540 18370 34620
rect 17690 34320 17730 34360
rect 17870 34320 17910 34360
rect 18040 34320 18080 34360
rect 18630 34320 18670 34360
rect 18810 34320 18850 34360
rect 18980 34320 19020 34360
rect 19750 34750 19810 34810
rect 20920 34900 20980 34960
rect 21190 34910 21230 34950
rect 19880 34770 19920 34810
rect 20020 34770 20060 34810
rect 19770 34620 19810 34660
rect 19580 34350 19640 34430
rect 20760 34450 20820 34530
rect 22540 35450 22580 35490
rect 22680 35450 22720 35490
rect 23000 35450 23040 35490
rect 22610 35320 22650 35360
rect 22200 35240 22270 35310
rect 23480 35450 23520 35490
rect 23620 35450 23660 35490
rect 23940 35450 23980 35490
rect 23550 35320 23590 35360
rect 22830 35160 22870 35200
rect 22430 34860 22470 34900
rect 23520 35170 23590 35240
rect 23370 34860 23410 34900
rect 23660 34860 23700 34900
rect 24730 35450 24770 35490
rect 24980 35480 25020 35520
rect 24090 34910 24130 34950
rect 24280 34910 24320 34950
rect 24480 34910 24520 34950
rect 25170 35330 25210 35370
rect 23240 34470 23300 34550
rect 22650 34320 22690 34360
rect 22830 34320 22870 34360
rect 23000 34320 23040 34360
rect 23590 34320 23630 34360
rect 23770 34320 23810 34360
rect 23940 34320 23980 34360
rect 24710 34750 24770 34810
rect 24840 34770 24880 34810
rect 24980 34770 25020 34810
rect 24730 34620 24770 34660
rect 24950 34300 25010 34380
rect 16510 34130 16570 34200
rect 16610 34130 16670 34200
rect 16710 34130 16770 34200
rect 16810 34130 16870 34200
rect 16910 34130 16970 34200
rect 17010 34130 17070 34200
rect 17110 34130 17170 34200
rect 17210 34130 17270 34200
rect 17310 34130 17370 34200
rect 17410 34130 17470 34200
rect 17510 34130 17570 34200
rect 17610 34130 17670 34200
rect 17710 34130 17770 34200
rect 17810 34130 17870 34200
rect 17910 34130 17970 34200
rect 18010 34130 18070 34200
rect 18110 34130 18170 34200
rect 18210 34130 18270 34200
rect 18310 34130 18370 34200
rect 18410 34130 18470 34200
rect 18510 34130 18570 34200
rect 18610 34130 18670 34200
rect 18710 34130 18770 34200
rect 18810 34130 18870 34200
rect 18910 34130 18970 34200
rect 19010 34130 19070 34200
rect 19110 34130 19170 34200
rect 19210 34130 19270 34200
rect 19310 34130 19370 34200
rect 19410 34130 19470 34200
rect 19510 34130 19570 34200
rect 19610 34130 19670 34200
rect 19710 34130 19770 34200
rect 19810 34130 19870 34200
rect 19910 34130 19970 34200
rect 20010 34130 20070 34200
rect 20110 34130 20170 34200
rect 20210 34130 20270 34200
rect 20310 34130 20370 34200
rect 20410 34130 20470 34200
rect 20510 34130 20570 34200
rect 20610 34130 20670 34200
rect 20710 34130 20770 34200
rect 20810 34130 20870 34200
rect 20910 34130 20970 34200
rect 21010 34130 21070 34200
rect 21110 34130 21170 34200
rect 21210 34130 21270 34200
rect 21310 34130 21370 34200
rect 21410 34130 21470 34200
rect 21510 34130 21570 34200
rect 21610 34130 21670 34200
rect 21710 34130 21770 34200
rect 21810 34130 21870 34200
rect 21910 34130 21970 34200
rect 22010 34130 22070 34200
rect 22110 34130 22170 34200
rect 22210 34130 22270 34200
rect 22310 34130 22370 34200
rect 22410 34130 22470 34200
rect 22510 34130 22570 34200
rect 22610 34130 22670 34200
rect 22710 34130 22770 34200
rect 22810 34130 22870 34200
rect 22910 34130 22970 34200
rect 23010 34130 23070 34200
rect 23110 34130 23170 34200
rect 23210 34130 23270 34200
rect 23310 34130 23370 34200
rect 23410 34130 23470 34200
rect 23510 34130 23570 34200
rect 23620 34130 23680 34200
rect 23720 34130 23780 34200
rect 23820 34130 23880 34200
rect 23920 34130 23980 34200
rect 24020 34130 24080 34200
rect 24120 34130 24180 34200
rect 24220 34130 24280 34200
rect 24320 34130 24380 34200
rect 24420 34130 24480 34200
rect 24520 34130 24580 34200
rect 24620 34130 24680 34200
rect 24720 34130 24780 34200
rect 24820 34130 24880 34200
rect 24920 34130 24980 34200
rect 25020 34130 25080 34200
rect 25120 34130 25180 34200
rect 25220 34130 25280 34200
rect 25320 34130 25380 34200
rect 6380 33980 6440 34040
rect 6480 33980 6540 34040
rect 6580 33980 6640 34040
rect 6680 33980 6740 34040
rect 6780 33980 6840 34040
rect 6880 33980 6940 34040
rect 6980 33980 7040 34040
rect 7080 33980 7140 34040
rect 7180 33980 7240 34040
rect 7280 33980 7340 34040
rect 7380 33980 7440 34040
rect 7480 33980 7540 34040
rect 7580 33980 7640 34040
rect 7680 33980 7740 34040
rect 7780 33980 7840 34040
rect 7880 33980 7940 34040
rect 7980 33980 8040 34040
rect 8080 33980 8140 34040
rect 8180 33980 8240 34040
rect 8280 33980 8340 34040
rect 8380 33980 8440 34040
rect 8480 33980 8540 34040
rect 8580 33980 8640 34040
rect 8680 33980 8740 34040
rect 8780 33980 8840 34040
rect 8880 33980 8940 34040
rect 8980 33980 9040 34040
rect 9080 33980 9140 34040
rect 9180 33980 9240 34040
rect 9280 33980 9340 34040
rect 9380 33980 9440 34040
rect 9480 33980 9540 34040
rect 9580 33980 9640 34040
rect 9680 33980 9740 34040
rect 9780 33980 9840 34040
rect 9880 33980 9940 34040
rect 9980 33980 10040 34040
rect 10080 33980 10140 34040
rect 10180 33980 10240 34040
rect 10280 33980 10340 34040
rect 10380 33980 10440 34040
rect 10480 33980 10540 34040
rect 10580 33980 10640 34040
rect 10680 33980 10740 34040
rect 10780 33980 10840 34040
rect 3810 33560 3870 33620
rect 3910 33560 3970 33620
rect 4010 33560 4070 33620
rect 4110 33560 4170 33620
rect 4210 33560 4270 33620
rect 4310 33560 4370 33620
rect 4410 33560 4470 33620
rect 4510 33560 4570 33620
rect 4610 33560 4670 33620
rect 4710 33560 4770 33620
rect 4810 33560 4870 33620
rect 4910 33560 4970 33620
rect 5010 33560 5070 33620
rect 5110 33560 5170 33620
rect 5210 33560 5270 33620
rect 5310 33560 5370 33620
rect 5410 33560 5470 33620
rect 5510 33560 5570 33620
rect 5610 33560 5670 33620
rect 5710 33560 5770 33620
rect 5810 33560 5870 33620
rect 5910 33560 5970 33620
rect 6010 33560 6070 33620
rect 6110 33560 6170 33620
rect 13768 32420 13848 32460
rect 14118 32340 14158 32380
rect 15650 32250 15710 32310
rect 14008 31900 14048 31940
rect 16120 32110 16180 32180
rect 16220 32110 16280 32180
rect 16320 32110 16380 32180
rect 16420 32110 16480 32180
rect 16520 32110 16580 32180
rect 16620 32110 16680 32180
rect 16720 32110 16780 32180
rect 16820 32110 16880 32180
rect 16920 32110 16980 32180
rect 17020 32110 17080 32180
rect 17120 32110 17180 32180
rect 17220 32110 17280 32180
rect 17320 32110 17380 32180
rect 17420 32110 17480 32180
rect 17520 32110 17580 32180
rect 17620 32110 17680 32180
rect 17720 32110 17780 32180
rect 17820 32110 17880 32180
rect 17920 32110 17980 32180
rect 18020 32110 18080 32180
rect 18120 32110 18180 32180
rect 18220 32110 18280 32180
rect 18320 32110 18380 32180
rect 18420 32110 18480 32180
rect 18520 32110 18580 32180
rect 18620 32110 18680 32180
rect 18720 32110 18780 32180
rect 18820 32110 18880 32180
rect 18920 32110 18980 32180
rect 19020 32110 19080 32180
rect 19120 32110 19180 32180
rect 19220 32110 19280 32180
rect 19320 32110 19380 32180
rect 19420 32110 19480 32180
rect 19520 32110 19580 32180
rect 19620 32110 19680 32180
rect 19720 32110 19780 32180
rect 19820 32110 19880 32180
rect 19920 32110 19980 32180
rect 20020 32110 20080 32180
rect 20120 32110 20180 32180
rect 20220 32110 20280 32180
rect 20320 32110 20380 32180
rect 20420 32110 20480 32180
rect 20520 32110 20580 32180
rect 20620 32110 20680 32180
rect 20720 32110 20780 32180
rect 20820 32110 20880 32180
rect 20920 32110 20980 32180
rect 21020 32110 21080 32180
rect 21120 32110 21180 32180
rect 21220 32110 21280 32180
rect 21320 32110 21380 32180
rect 21420 32110 21480 32180
rect 21520 32110 21580 32180
rect 21620 32110 21680 32180
rect 21720 32110 21780 32180
rect 21820 32110 21880 32180
rect 21920 32110 21980 32180
rect 22020 32110 22080 32180
rect 22120 32110 22180 32180
rect 22220 32110 22280 32180
rect 22320 32110 22380 32180
rect 22420 32110 22480 32180
rect 22520 32110 22580 32180
rect 22620 32110 22680 32180
rect 22720 32110 22780 32180
rect 22820 32110 22880 32180
rect 22920 32110 22980 32180
rect 23020 32110 23080 32180
rect 23120 32110 23180 32180
rect 23220 32110 23280 32180
rect 23320 32110 23380 32180
rect 23420 32110 23480 32180
rect 23520 32110 23580 32180
rect 23620 32110 23680 32180
rect 23720 32110 23780 32180
rect 23820 32110 23880 32180
rect 23920 32110 23980 32180
rect 24020 32110 24080 32180
rect 24120 32110 24180 32180
rect 24220 32110 24280 32180
rect 24320 32110 24380 32180
rect 24420 32110 24480 32180
rect 24520 32110 24580 32180
rect 24620 32110 24680 32180
rect 24720 32110 24780 32180
rect 24820 32110 24880 32180
rect 24920 32110 24980 32180
rect 25020 32110 25080 32180
rect 25120 32110 25180 32180
rect 25220 32110 25280 32180
rect 25320 32110 25380 32180
rect 14400 31950 14510 32010
rect 15590 31940 15650 32020
rect 14228 31850 14268 31890
rect 14118 31750 14158 31790
rect 2210 31670 2270 31730
rect 2310 31670 2370 31730
rect 2410 31670 2470 31730
rect 2510 31670 2570 31730
rect 2610 31670 2670 31730
rect 2710 31670 2770 31730
rect 2810 31670 2870 31730
rect 2910 31670 2970 31730
rect 3010 31670 3070 31730
rect 3110 31670 3170 31730
rect 3210 31670 3270 31730
rect 3310 31670 3370 31730
rect 3410 31670 3470 31730
rect 3510 31670 3570 31730
rect 3610 31670 3670 31730
rect 3710 31670 3770 31730
rect 3810 31670 3870 31730
rect 3910 31670 3970 31730
rect 4010 31670 4070 31730
rect 4110 31670 4170 31730
rect 4210 31670 4270 31730
rect 4310 31670 4370 31730
rect 4410 31670 4470 31730
rect 4510 31670 4570 31730
rect 4610 31670 4670 31730
rect 4710 31670 4770 31730
rect 4810 31670 4870 31730
rect 4910 31670 4970 31730
rect 5010 31670 5070 31730
rect 5110 31670 5170 31730
rect 5210 31670 5270 31730
rect 5310 31670 5370 31730
rect 5410 31670 5470 31730
rect 5510 31670 5570 31730
rect 5610 31670 5670 31730
rect 5710 31670 5770 31730
rect 5810 31670 5870 31730
rect 5910 31670 5970 31730
rect 6010 31670 6070 31730
rect 6110 31670 6170 31730
rect 6210 31670 6270 31730
rect 2160 30690 2210 30740
rect 2960 30680 3020 30740
rect 6470 31320 6530 31380
rect 6580 31320 6640 31380
rect 6690 31320 6750 31380
rect 6800 31320 6860 31380
rect 6910 31320 6970 31380
rect 7020 31320 7080 31380
rect 7130 31320 7190 31380
rect 7240 31320 7300 31380
rect 7350 31320 7410 31380
rect 7460 31320 7520 31380
rect 7570 31320 7630 31380
rect 7680 31320 7740 31380
rect 7790 31320 7850 31380
rect 7900 31320 7960 31380
rect 8010 31320 8070 31380
rect 8120 31320 8180 31380
rect 8230 31320 8290 31380
rect 8340 31320 8400 31380
rect 8450 31320 8510 31380
rect 8560 31320 8620 31380
rect 8670 31320 8730 31380
rect 8780 31320 8840 31380
rect 8890 31320 8950 31380
rect 9000 31320 9060 31380
rect 9110 31320 9170 31380
rect 9220 31320 9280 31380
rect 9330 31320 9390 31380
rect 9440 31320 9500 31380
rect 9550 31320 9610 31380
rect 9660 31320 9720 31380
rect 9770 31320 9830 31380
rect 9880 31320 9940 31380
rect 9990 31320 10050 31380
rect 10100 31320 10160 31380
rect 10210 31320 10270 31380
rect 10320 31320 10380 31380
rect 10430 31320 10490 31380
rect 10540 31320 10600 31380
rect 10650 31320 10710 31380
rect 10760 31320 10820 31380
rect 10880 31320 10940 31380
rect 10990 31320 11050 31380
rect 11100 31320 11160 31380
rect 16450 31390 16510 31450
rect 17140 31390 17180 31430
rect 6310 30660 6360 30710
rect 6400 30660 6440 30700
rect 9120 30760 9160 30800
rect 14118 31270 14158 31310
rect 6700 30660 6740 30700
rect 6780 30660 6820 30700
rect 3730 30560 3770 30600
rect 3820 30560 3860 30600
rect 4590 30560 4640 30610
rect 4680 30560 4730 30610
rect 5450 30560 5500 30610
rect 5540 30560 5590 30610
rect 7280 30650 7320 30690
rect 7360 30650 7400 30690
rect 7660 30650 7700 30690
rect 7740 30650 7780 30690
rect 8040 30650 8080 30690
rect 8120 30650 8160 30690
rect 8420 30650 8460 30690
rect 8500 30650 8540 30690
rect 8750 30650 8790 30690
rect 8860 30650 8900 30690
rect 7240 30000 7280 30040
rect 9360 30650 9400 30690
rect 9440 30650 9480 30690
rect 9740 30650 9780 30690
rect 9820 30650 9860 30690
rect 10120 30650 10160 30690
rect 10200 30650 10240 30690
rect 10500 30650 10540 30690
rect 10580 30650 10620 30690
rect 10880 30650 10920 30690
rect 10960 30650 11000 30690
rect 11240 30660 11300 30720
rect 15400 30210 15470 30280
rect 17240 31230 17310 31300
rect 17580 31390 17620 31430
rect 17720 31390 17760 31430
rect 18040 31390 18080 31430
rect 17650 31260 17690 31300
rect 18520 31390 18560 31430
rect 18660 31390 18700 31430
rect 18980 31390 19020 31430
rect 18590 31260 18630 31300
rect 17870 31100 17910 31140
rect 17470 30800 17510 30840
rect 18540 31080 18610 31150
rect 18410 30800 18450 30840
rect 18700 30800 18740 30840
rect 20030 31390 20070 31430
rect 20280 31400 20320 31440
rect 19130 30850 19170 30890
rect 19320 30850 19360 30890
rect 19460 30850 19500 30890
rect 19580 30850 19620 30890
rect 19780 30850 19820 30890
rect 20470 31200 20510 31240
rect 21490 31380 21530 31420
rect 22160 31380 22200 31420
rect 18240 30400 18310 30480
rect 17690 30260 17730 30300
rect 17870 30260 17910 30300
rect 18040 30260 18080 30300
rect 18630 30260 18670 30300
rect 18810 30260 18850 30300
rect 18980 30260 19020 30300
rect 20010 30690 20070 30750
rect 20980 30840 21040 30900
rect 20140 30710 20180 30750
rect 20280 30710 20320 30750
rect 20030 30560 20070 30600
rect 20740 30760 20800 30840
rect 21250 30850 21290 30890
rect 20560 30380 20620 30460
rect 20740 30380 20800 30460
rect 22260 31230 22330 31300
rect 22600 31380 22640 31420
rect 22740 31380 22780 31420
rect 23060 31380 23100 31420
rect 22670 31250 22710 31290
rect 23540 31380 23580 31420
rect 23680 31380 23720 31420
rect 24000 31380 24040 31420
rect 23610 31250 23650 31290
rect 22890 31090 22930 31130
rect 22490 30790 22530 30830
rect 23570 31080 23640 31150
rect 23430 30790 23470 30830
rect 23720 30790 23760 30830
rect 24990 31380 25030 31420
rect 25240 31410 25280 31450
rect 24150 30840 24190 30880
rect 24340 30840 24380 30880
rect 24490 30840 24530 30880
rect 24600 30840 24640 30880
rect 24740 30840 24780 30880
rect 25430 31260 25470 31300
rect 23260 30400 23320 30480
rect 22710 30250 22750 30290
rect 22890 30250 22930 30290
rect 23060 30250 23100 30290
rect 23650 30250 23690 30290
rect 23830 30250 23870 30290
rect 24000 30250 24040 30290
rect 24970 30680 25030 30740
rect 25100 30700 25140 30740
rect 25240 30700 25280 30740
rect 24990 30550 25030 30590
rect 14870 30060 14930 30130
rect 14970 30060 15030 30130
rect 15070 30060 15130 30130
rect 15170 30060 15230 30130
rect 15270 30060 15330 30130
rect 15370 30060 15430 30130
rect 15470 30060 15530 30130
rect 15570 30060 15630 30130
rect 15670 30060 15730 30130
rect 15780 30060 15840 30130
rect 15880 30060 15940 30130
rect 15990 30060 16050 30130
rect 16130 30060 16190 30130
rect 16270 30060 16330 30130
rect 16370 30060 16430 30130
rect 16470 30060 16530 30130
rect 16570 30060 16630 30130
rect 16670 30060 16730 30130
rect 16770 30060 16830 30130
rect 16870 30060 16930 30130
rect 16970 30060 17030 30130
rect 17070 30060 17130 30130
rect 17170 30060 17230 30130
rect 17270 30060 17330 30130
rect 17370 30060 17430 30130
rect 17470 30060 17530 30130
rect 17570 30060 17630 30130
rect 17670 30060 17730 30130
rect 17770 30060 17830 30130
rect 17870 30060 17930 30130
rect 17970 30060 18030 30130
rect 18070 30060 18130 30130
rect 18170 30060 18230 30130
rect 18270 30060 18330 30130
rect 18370 30060 18430 30130
rect 18470 30060 18530 30130
rect 18570 30060 18630 30130
rect 18670 30060 18730 30130
rect 18770 30060 18830 30130
rect 18870 30060 18930 30130
rect 18970 30060 19030 30130
rect 19070 30060 19130 30130
rect 19170 30060 19230 30130
rect 19270 30060 19330 30130
rect 19370 30060 19430 30130
rect 19470 30060 19530 30130
rect 19570 30060 19630 30130
rect 19670 30060 19730 30130
rect 19770 30060 19830 30130
rect 19870 30060 19930 30130
rect 19970 30060 20030 30130
rect 20070 30060 20130 30130
rect 20170 30060 20230 30130
rect 20270 30060 20330 30130
rect 20370 30060 20430 30130
rect 20470 30060 20530 30130
rect 20570 30060 20630 30130
rect 20670 30060 20730 30130
rect 20770 30060 20830 30130
rect 20870 30060 20930 30130
rect 20970 30060 21030 30130
rect 21070 30060 21130 30130
rect 21170 30060 21230 30130
rect 21270 30060 21330 30130
rect 21370 30060 21430 30130
rect 21470 30060 21530 30130
rect 21570 30060 21630 30130
rect 21670 30060 21730 30130
rect 21770 30060 21830 30130
rect 21870 30060 21930 30130
rect 21970 30060 22030 30130
rect 22070 30060 22130 30130
rect 22170 30060 22230 30130
rect 22270 30060 22330 30130
rect 22370 30060 22430 30130
rect 22470 30060 22530 30130
rect 22570 30060 22630 30130
rect 22670 30060 22730 30130
rect 22770 30060 22830 30130
rect 22870 30060 22930 30130
rect 22970 30060 23030 30130
rect 23070 30060 23130 30130
rect 23170 30060 23230 30130
rect 23270 30060 23330 30130
rect 23370 30060 23430 30130
rect 23470 30060 23530 30130
rect 23570 30060 23630 30130
rect 23670 30060 23730 30130
rect 23770 30060 23830 30130
rect 23870 30060 23930 30130
rect 23970 30060 24030 30130
rect 24070 30060 24130 30130
rect 24170 30060 24230 30130
rect 24270 30060 24330 30130
rect 24370 30060 24430 30130
rect 24470 30060 24530 30130
rect 24570 30060 24630 30130
rect 24670 30060 24730 30130
rect 24770 30060 24830 30130
rect 24870 30060 24930 30130
rect 24970 30060 25030 30130
rect 25070 30060 25130 30130
rect 25170 30060 25230 30130
rect 25270 30060 25330 30130
rect 25370 30060 25430 30130
rect 25470 30060 25530 30130
rect 25570 30060 25630 30130
rect 6440 29840 6500 29900
rect 6540 29840 6600 29900
rect 6640 29840 6700 29900
rect 6740 29840 6800 29900
rect 6840 29840 6900 29900
rect 6940 29840 7000 29900
rect 7040 29840 7100 29900
rect 7140 29840 7200 29900
rect 7240 29840 7300 29900
rect 7340 29840 7400 29900
rect 7440 29840 7500 29900
rect 7540 29840 7600 29900
rect 7640 29840 7700 29900
rect 7740 29840 7800 29900
rect 7840 29840 7900 29900
rect 7940 29840 8000 29900
rect 8040 29840 8100 29900
rect 8140 29840 8200 29900
rect 8240 29840 8300 29900
rect 8340 29840 8400 29900
rect 8440 29840 8500 29900
rect 8540 29840 8600 29900
rect 8640 29840 8700 29900
rect 8740 29840 8800 29900
rect 8840 29840 8900 29900
rect 8940 29840 9000 29900
rect 9040 29840 9100 29900
rect 9140 29840 9200 29900
rect 9240 29840 9300 29900
rect 9340 29840 9400 29900
rect 9440 29840 9500 29900
rect 9540 29840 9600 29900
rect 9640 29840 9700 29900
rect 9740 29840 9800 29900
rect 9840 29840 9900 29900
rect 9940 29840 10000 29900
rect 10040 29840 10100 29900
rect 10140 29840 10200 29900
rect 10240 29840 10300 29900
rect 10340 29840 10400 29900
rect 10440 29840 10500 29900
rect 10540 29840 10600 29900
rect 10640 29840 10700 29900
rect 10740 29840 10800 29900
rect 10840 29840 10900 29900
rect 10940 29840 11000 29900
rect 11040 29840 11100 29900
rect 11140 29840 11200 29900
rect 2210 29310 2270 29370
rect 2310 29310 2370 29370
rect 2410 29310 2470 29370
rect 2510 29310 2570 29370
rect 2610 29310 2670 29370
rect 2710 29310 2770 29370
rect 2810 29310 2870 29370
rect 2910 29310 2970 29370
rect 3010 29310 3070 29370
rect 3110 29310 3170 29370
rect 3210 29310 3270 29370
rect 3310 29310 3370 29370
rect 3410 29310 3470 29370
rect 3510 29310 3570 29370
rect 3610 29310 3670 29370
rect 3710 29310 3770 29370
rect 3810 29310 3870 29370
rect 3910 29310 3970 29370
rect 4010 29310 4070 29370
rect 4110 29310 4170 29370
rect 4210 29310 4270 29370
rect 4310 29310 4370 29370
rect 4410 29310 4470 29370
rect 4510 29310 4570 29370
rect 4610 29310 4670 29370
rect 4710 29310 4770 29370
rect 4810 29310 4870 29370
rect 4910 29310 4970 29370
rect 5010 29310 5070 29370
rect 5110 29310 5170 29370
rect 5210 29310 5270 29370
rect 5310 29310 5370 29370
rect 5410 29310 5470 29370
rect 5510 29310 5570 29370
rect 5610 29310 5670 29370
rect 5710 29310 5770 29370
rect 5810 29310 5870 29370
rect 5910 29310 5970 29370
rect 6010 29310 6070 29370
rect 6110 29310 6170 29370
rect 6210 29310 6270 29370
rect 7360 26570 7400 26610
rect 7440 26570 7480 26610
rect 7520 26570 7560 26610
rect 7600 26570 7640 26610
rect 7680 26570 7720 26610
rect 7760 26570 7800 26610
rect 7840 26570 7880 26610
rect 7920 26570 7960 26610
rect 8000 26570 8040 26610
rect 8080 26570 8120 26610
rect 8160 26570 8200 26610
rect 8240 26570 8280 26610
rect 8320 26570 8360 26610
rect 8400 26570 8440 26610
rect 8480 26570 8520 26610
rect 8560 26570 8600 26610
rect 8640 26570 8680 26610
rect 8720 26570 8760 26610
rect 8800 26570 8840 26610
rect 8880 26570 8920 26610
rect 8960 26570 9000 26610
rect 9040 26570 9080 26610
rect 9120 26570 9160 26610
rect 9200 26570 9240 26610
rect 9280 26570 9320 26610
rect 9360 26570 9400 26610
rect 9440 26570 9480 26610
rect 9520 26570 9560 26610
rect 9600 26570 9640 26610
rect 9680 26570 9720 26610
rect 9760 26570 9800 26610
rect 9840 26570 9880 26610
rect 9920 26570 9960 26610
rect 10000 26570 10040 26610
rect 10080 26570 10120 26610
rect 10160 26570 10200 26610
rect 10240 26570 10280 26610
rect 10320 26570 10360 26610
rect 10400 26570 10440 26610
rect 10480 26570 10520 26610
rect 10560 26570 10600 26610
rect 10640 26570 10680 26610
rect 10720 26570 10760 26610
rect 10800 26570 10840 26610
rect 10880 26570 10920 26610
rect 10960 26570 11000 26610
rect 11040 26570 11080 26610
rect 11120 26570 11160 26610
rect 11200 26570 11240 26610
rect 11280 26570 11320 26610
rect 11360 26570 11400 26610
rect 11440 26570 11480 26610
rect 11520 26570 11560 26610
rect 11600 26570 11640 26610
rect 11680 26570 11720 26610
rect 11760 26570 11800 26610
rect 11840 26570 11880 26610
rect 11920 26570 11960 26610
rect 12000 26570 12040 26610
rect 12080 26570 12120 26610
rect 12160 26570 12200 26610
rect 12240 26570 12280 26610
rect 12320 26570 12360 26610
rect 12400 26570 12440 26610
rect 12480 26570 12520 26610
rect 12560 26570 12600 26610
rect 12640 26570 12680 26610
rect 12720 26570 12760 26610
rect 12800 26570 12840 26610
rect 12880 26570 12920 26610
rect 12960 26570 13000 26610
rect 13040 26570 13080 26610
rect 13120 26570 13160 26610
rect 13200 26570 13240 26610
rect 13280 26570 13320 26610
rect 13360 26570 13400 26610
rect 13440 26570 13480 26610
rect 13520 26570 13560 26610
rect 13600 26570 13640 26610
rect 13680 26570 13720 26610
rect 13760 26570 13800 26610
rect 13840 26570 13880 26610
rect 13920 26570 13960 26610
rect 14000 26570 14040 26610
rect 14080 26570 14120 26610
rect 14160 26570 14200 26610
rect 14240 26570 14280 26610
rect 14320 26570 14360 26610
rect 14400 26570 14440 26610
rect 14480 26570 14520 26610
rect 14560 26570 14600 26610
rect 14640 26570 14680 26610
rect 14720 26570 14760 26610
rect 14800 26570 14840 26610
rect 14880 26570 14920 26610
rect 14960 26570 15000 26610
rect 15040 26570 15080 26610
rect 15120 26570 15160 26610
rect 15200 26570 15240 26610
rect 15280 26570 15320 26610
rect 15360 26570 15400 26610
rect 15440 26570 15480 26610
rect 15520 26570 15560 26610
rect 15600 26570 15640 26610
rect 15680 26570 15720 26610
rect 15760 26570 15800 26610
rect 15840 26570 15880 26610
rect 15920 26570 15960 26610
rect 16000 26570 16040 26610
rect 16080 26570 16120 26610
rect 16160 26570 16200 26610
rect 16240 26570 16280 26610
rect 16320 26570 16360 26610
rect 16400 26570 16440 26610
rect 16480 26570 16520 26610
rect 16560 26570 16600 26610
rect 16640 26570 16680 26610
rect 16720 26570 16760 26610
rect 16800 26570 16840 26610
rect 16880 26570 16920 26610
rect 16960 26570 17000 26610
rect 17040 26570 17080 26610
rect 17120 26570 17160 26610
rect 17200 26570 17240 26610
rect 17280 26570 17320 26610
rect 17360 26570 17400 26610
rect 17440 26570 17480 26610
rect 17520 26570 17560 26610
rect 17600 26570 17640 26610
rect 17680 26570 17720 26610
rect 17760 26570 17800 26610
rect 17840 26570 17880 26610
rect 17920 26570 17960 26610
rect 18000 26570 18040 26610
rect 18080 26570 18120 26610
rect 18160 26570 18200 26610
rect 18240 26570 18280 26610
rect 18320 26570 18360 26610
rect 18400 26570 18440 26610
rect 18480 26570 18520 26610
rect 18560 26570 18600 26610
rect 18640 26570 18680 26610
rect 18720 26570 18760 26610
rect 18800 26570 18840 26610
rect 18880 26570 18920 26610
rect 18960 26570 19000 26610
rect 19040 26570 19080 26610
rect 19120 26570 19160 26610
rect 19200 26570 19240 26610
rect 19280 26570 19320 26610
rect 19360 26570 19400 26610
rect 19440 26570 19480 26610
rect 19520 26570 19560 26610
rect 19600 26570 19640 26610
rect 19680 26570 19720 26610
rect 19760 26570 19800 26610
rect 19840 26570 19880 26610
rect 19920 26570 19960 26610
rect 20000 26570 20040 26610
rect 20080 26570 20120 26610
rect 20160 26570 20200 26610
rect 20240 26570 20280 26610
rect 20320 26570 20360 26610
rect 20400 26570 20440 26610
rect 20480 26570 20520 26610
rect 20560 26570 20600 26610
rect 6300 25500 6360 25560
rect 7080 25500 7140 25560
rect 7290 25130 7350 25190
rect 7820 25500 7880 25560
rect 8500 24900 8540 24940
rect 8800 24900 8840 24940
rect 8880 24900 8920 24940
rect 8990 24890 9050 24950
rect 9220 24910 9260 24950
rect 8080 24800 8140 24870
rect 8650 24820 8690 24860
rect 7570 24710 7630 24770
rect 8200 24670 8260 24730
rect 9680 25910 9720 25950
rect 9680 25020 9720 25060
rect 9940 25910 9980 25950
rect 9940 25020 9980 25060
rect 10670 25910 10710 25950
rect 10670 25020 10710 25060
rect 10930 25910 10970 25950
rect 10930 25020 10970 25060
rect 11670 25910 11710 25950
rect 11670 25020 11710 25060
rect 11930 25910 11970 25950
rect 11930 25020 11970 25060
rect 9580 24900 9620 24940
rect 10080 24910 10120 24950
rect 10160 24910 10200 24950
rect 10460 24910 10500 24950
rect 10570 24900 10610 24940
rect 11070 24910 11110 24950
rect 11150 24910 11190 24950
rect 11450 24910 11490 24950
rect 11570 24900 11610 24940
rect 12070 24910 12110 24950
rect 12150 24910 12190 24950
rect 12450 24910 12490 24950
rect 12530 24910 12570 24950
rect 12820 24900 12860 24940
rect 12900 24900 12940 24940
rect 9840 24800 9880 24840
rect 9100 24560 9150 24610
rect 9090 24380 9160 24440
rect 10410 24790 10480 24850
rect 10830 24800 10870 24840
rect 11410 24790 11480 24850
rect 11830 24800 11870 24840
rect 13230 25890 13270 25930
rect 13230 25000 13270 25040
rect 13000 24900 13040 24940
rect 13130 24900 13170 24940
rect 13570 25890 13610 25930
rect 13790 25890 13830 25930
rect 13570 25000 13610 25040
rect 13790 25000 13830 25040
rect 13340 24900 13380 24940
rect 13470 24900 13510 24940
rect 14130 25910 14170 25950
rect 14350 25910 14390 25950
rect 14570 25910 14610 25950
rect 14790 25910 14830 25950
rect 14130 25020 14170 25060
rect 14350 25020 14390 25060
rect 14570 25020 14610 25060
rect 14790 25020 14830 25060
rect 13900 24900 13940 24940
rect 14030 24900 14070 24940
rect 15190 25910 15230 25950
rect 15410 25910 15450 25950
rect 15630 25910 15670 25950
rect 15850 25910 15890 25950
rect 16070 25910 16110 25950
rect 16290 25910 16330 25950
rect 16510 25910 16550 25950
rect 16730 25910 16770 25950
rect 15190 25020 15230 25060
rect 15410 25020 15450 25060
rect 15630 25020 15670 25060
rect 15850 25020 15890 25060
rect 16070 25020 16110 25060
rect 16290 25020 16330 25060
rect 16510 25020 16550 25060
rect 16730 25020 16770 25060
rect 14900 24900 14940 24940
rect 15090 24900 15130 24940
rect 17140 25910 17180 25950
rect 17360 25910 17400 25950
rect 17580 25910 17620 25950
rect 17800 25910 17840 25950
rect 18020 25910 18060 25950
rect 18240 25910 18280 25950
rect 18460 25910 18500 25950
rect 18680 25910 18720 25950
rect 18900 25910 18940 25950
rect 19120 25910 19160 25950
rect 19340 25910 19380 25950
rect 19560 25910 19600 25950
rect 19780 25910 19820 25950
rect 20000 25910 20040 25950
rect 20220 25910 20260 25950
rect 20440 25910 20480 25950
rect 17140 25020 17180 25060
rect 17360 25020 17400 25060
rect 17580 25020 17620 25060
rect 17800 25020 17840 25060
rect 18020 25020 18060 25060
rect 18240 25020 18280 25060
rect 18460 25020 18500 25060
rect 18680 25020 18720 25060
rect 18900 25020 18940 25060
rect 19120 25020 19160 25060
rect 19340 25020 19380 25060
rect 19560 25020 19600 25060
rect 19780 25020 19820 25060
rect 20000 25020 20040 25060
rect 20220 25020 20260 25060
rect 20440 25020 20480 25060
rect 16890 24890 16940 24940
rect 17040 24900 17080 24940
rect 20600 24890 20650 24940
rect 7320 24250 7360 24290
rect 7400 24250 7440 24290
rect 7480 24250 7520 24290
rect 7560 24250 7600 24290
rect 7640 24250 7680 24290
rect 7720 24250 7760 24290
rect 7800 24250 7840 24290
rect 7890 24250 7930 24290
rect 7970 24250 8010 24290
rect 8050 24250 8090 24290
rect 8130 24250 8170 24290
rect 8210 24250 8250 24290
rect 8290 24250 8330 24290
rect 8400 24250 8440 24290
rect 8520 24250 8560 24290
rect 8600 24250 8640 24290
rect 8680 24250 8720 24290
rect 8760 24250 8800 24290
rect 8840 24250 8880 24290
rect 8920 24250 8960 24290
rect 9000 24250 9040 24290
rect 9080 24250 9120 24290
rect 9160 24250 9200 24290
rect 9270 24250 9310 24290
rect 9350 24250 9390 24290
rect 9430 24250 9470 24290
rect 9510 24250 9550 24290
rect 9590 24250 9630 24290
rect 9670 24250 9710 24290
rect 9750 24250 9790 24290
rect 9830 24250 9870 24290
rect 9910 24250 9950 24290
rect 9990 24250 10030 24290
rect 10070 24250 10110 24290
rect 10150 24250 10190 24290
rect 10230 24250 10270 24290
rect 10310 24250 10350 24290
rect 10390 24250 10430 24290
rect 10470 24250 10510 24290
rect 10550 24250 10590 24290
rect 10630 24250 10670 24290
rect 10710 24250 10750 24290
rect 10790 24250 10830 24290
rect 10870 24250 10910 24290
rect 10950 24250 10990 24290
rect 11030 24250 11070 24290
rect 11110 24250 11150 24290
rect 11190 24250 11230 24290
rect 11270 24250 11310 24290
rect 11350 24250 11390 24290
rect 11430 24250 11470 24290
rect 11510 24250 11550 24290
rect 11590 24250 11630 24290
rect 11670 24250 11710 24290
rect 11750 24250 11790 24290
rect 11830 24250 11870 24290
rect 11910 24250 11950 24290
rect 11990 24250 12030 24290
rect 12070 24250 12110 24290
rect 12150 24250 12190 24290
rect 12230 24250 12270 24290
rect 12310 24250 12350 24290
rect 12390 24250 12430 24290
rect 12470 24250 12510 24290
rect 12550 24250 12590 24290
rect 12630 24250 12670 24290
rect 12710 24250 12750 24290
rect 12790 24250 12830 24290
rect 12870 24250 12910 24290
rect 12950 24250 12990 24290
rect 13030 24250 13070 24290
rect 13110 24250 13150 24290
rect 13190 24250 13230 24290
rect 13270 24250 13310 24290
rect 13350 24250 13390 24290
rect 13430 24250 13470 24290
rect 13510 24250 13550 24290
rect 13590 24250 13630 24290
rect 13670 24250 13710 24290
rect 13750 24250 13790 24290
rect 13830 24250 13870 24290
rect 13910 24250 13950 24290
rect 13990 24250 14030 24290
rect 14070 24250 14110 24290
rect 14150 24250 14190 24290
rect 14230 24250 14270 24290
rect 14310 24250 14350 24290
rect 14390 24250 14430 24290
rect 14470 24250 14510 24290
rect 14550 24250 14590 24290
rect 14630 24250 14670 24290
rect 14710 24250 14750 24290
rect 14790 24250 14830 24290
rect 14870 24250 14910 24290
rect 14950 24250 14990 24290
rect 15030 24250 15070 24290
rect 15110 24250 15150 24290
rect 15190 24250 15230 24290
rect 15270 24250 15310 24290
rect 15350 24250 15390 24290
rect 15430 24250 15470 24290
rect 15510 24250 15550 24290
rect 15590 24250 15630 24290
rect 15670 24250 15710 24290
rect 15750 24250 15790 24290
rect 15830 24250 15870 24290
rect 15910 24250 15950 24290
rect 15990 24250 16030 24290
rect 16070 24250 16110 24290
rect 16150 24250 16190 24290
rect 16230 24250 16270 24290
rect 16310 24250 16350 24290
rect 16390 24250 16430 24290
rect 16470 24250 16510 24290
rect 16550 24250 16590 24290
rect 16630 24250 16670 24290
rect 16710 24250 16750 24290
rect 16790 24250 16830 24290
rect 16870 24250 16910 24290
rect 16950 24250 16990 24290
rect 17030 24250 17070 24290
rect 17110 24250 17150 24290
rect 17190 24250 17230 24290
rect 17270 24250 17310 24290
rect 17350 24250 17390 24290
rect 17430 24250 17470 24290
rect 17510 24250 17550 24290
rect 17590 24250 17630 24290
rect 17670 24250 17710 24290
rect 17750 24250 17790 24290
rect 17830 24250 17870 24290
rect 17910 24250 17950 24290
rect 17990 24250 18030 24290
rect 18070 24250 18110 24290
rect 18150 24250 18190 24290
rect 18230 24250 18270 24290
rect 18310 24250 18350 24290
rect 18390 24250 18430 24290
rect 18470 24250 18510 24290
rect 18550 24250 18590 24290
rect 18630 24250 18670 24290
rect 18710 24250 18750 24290
rect 18790 24250 18830 24290
rect 18870 24250 18910 24290
rect 18950 24250 18990 24290
rect 19030 24250 19070 24290
rect 19110 24250 19150 24290
rect 19190 24250 19230 24290
rect 19270 24250 19310 24290
rect 19350 24250 19390 24290
rect 19430 24250 19470 24290
rect 19510 24250 19550 24290
rect 19590 24250 19630 24290
rect 19670 24250 19710 24290
rect 19750 24250 19790 24290
rect 19830 24250 19870 24290
rect 19910 24250 19950 24290
rect 19990 24250 20030 24290
rect 20070 24250 20110 24290
rect 20150 24250 20190 24290
rect 20230 24250 20270 24290
rect 20310 24250 20350 24290
rect 20390 24250 20430 24290
rect 20470 24250 20510 24290
rect 20550 24250 20590 24290
rect 7310 23280 7350 23320
rect 7390 23280 7430 23320
rect 7470 23280 7510 23320
rect 7550 23280 7590 23320
rect 7630 23280 7670 23320
rect 7710 23280 7750 23320
rect 7790 23280 7830 23320
rect 7870 23280 7910 23320
rect 7950 23280 7990 23320
rect 8030 23280 8070 23320
rect 8110 23280 8150 23320
rect 8190 23280 8230 23320
rect 8270 23280 8310 23320
rect 8350 23280 8390 23320
rect 8430 23280 8470 23320
rect 8520 23280 8560 23320
rect 8600 23280 8640 23320
rect 8680 23280 8720 23320
rect 8760 23280 8800 23320
rect 8840 23280 8880 23320
rect 8920 23280 8960 23320
rect 9000 23280 9040 23320
rect 9080 23280 9120 23320
rect 9160 23280 9200 23320
rect 9270 23280 9310 23320
rect 9350 23280 9390 23320
rect 9430 23280 9470 23320
rect 9510 23280 9550 23320
rect 9590 23280 9630 23320
rect 9670 23280 9710 23320
rect 9750 23280 9790 23320
rect 9830 23280 9870 23320
rect 9910 23280 9950 23320
rect 9990 23280 10030 23320
rect 10070 23280 10110 23320
rect 10150 23280 10190 23320
rect 10230 23280 10270 23320
rect 10310 23280 10350 23320
rect 10390 23280 10430 23320
rect 10470 23280 10510 23320
rect 10550 23280 10590 23320
rect 10630 23280 10670 23320
rect 10710 23280 10750 23320
rect 10790 23280 10830 23320
rect 10870 23280 10910 23320
rect 10950 23280 10990 23320
rect 11030 23280 11070 23320
rect 11110 23280 11150 23320
rect 11190 23280 11230 23320
rect 11270 23280 11310 23320
rect 11350 23280 11390 23320
rect 11430 23280 11470 23320
rect 11510 23280 11550 23320
rect 11590 23280 11630 23320
rect 11670 23280 11710 23320
rect 11750 23280 11790 23320
rect 11830 23280 11870 23320
rect 11910 23280 11950 23320
rect 11990 23280 12030 23320
rect 12070 23280 12110 23320
rect 12150 23280 12190 23320
rect 12230 23280 12270 23320
rect 12310 23280 12350 23320
rect 12390 23280 12430 23320
rect 12470 23280 12510 23320
rect 12550 23280 12590 23320
rect 12630 23280 12670 23320
rect 12710 23280 12750 23320
rect 12790 23280 12830 23320
rect 12870 23280 12910 23320
rect 12950 23280 12990 23320
rect 13030 23280 13070 23320
rect 13110 23280 13150 23320
rect 13190 23280 13230 23320
rect 13270 23280 13310 23320
rect 13350 23280 13390 23320
rect 13430 23280 13470 23320
rect 13510 23280 13550 23320
rect 13590 23280 13630 23320
rect 13670 23280 13710 23320
rect 13750 23280 13790 23320
rect 13830 23280 13870 23320
rect 13910 23280 13950 23320
rect 13990 23280 14030 23320
rect 14070 23280 14110 23320
rect 14150 23280 14190 23320
rect 14230 23280 14270 23320
rect 14310 23280 14350 23320
rect 14390 23280 14430 23320
rect 14470 23280 14510 23320
rect 14550 23280 14590 23320
rect 14630 23280 14670 23320
rect 14710 23280 14750 23320
rect 14790 23280 14830 23320
rect 14870 23280 14910 23320
rect 14950 23280 14990 23320
rect 15030 23280 15070 23320
rect 15110 23280 15150 23320
rect 15190 23280 15230 23320
rect 15270 23280 15310 23320
rect 15350 23280 15390 23320
rect 15430 23280 15470 23320
rect 15510 23280 15550 23320
rect 15590 23280 15630 23320
rect 15670 23280 15710 23320
rect 15750 23280 15790 23320
rect 15830 23280 15870 23320
rect 15910 23280 15950 23320
rect 15990 23280 16030 23320
rect 16070 23280 16110 23320
rect 16150 23280 16190 23320
rect 16230 23280 16270 23320
rect 16310 23280 16350 23320
rect 16390 23280 16430 23320
rect 16470 23280 16510 23320
rect 16550 23280 16590 23320
rect 16630 23280 16670 23320
rect 16710 23280 16750 23320
rect 16790 23280 16830 23320
rect 16870 23280 16910 23320
rect 16950 23280 16990 23320
rect 17030 23280 17070 23320
rect 17110 23280 17150 23320
rect 17190 23280 17230 23320
rect 17270 23280 17310 23320
rect 17350 23280 17390 23320
rect 17430 23280 17470 23320
rect 17510 23280 17550 23320
rect 17590 23280 17630 23320
rect 17670 23280 17710 23320
rect 17750 23280 17790 23320
rect 17830 23280 17870 23320
rect 17910 23280 17950 23320
rect 17990 23280 18030 23320
rect 18070 23280 18110 23320
rect 18150 23280 18190 23320
rect 18230 23280 18270 23320
rect 18310 23280 18350 23320
rect 18390 23280 18430 23320
rect 18470 23280 18510 23320
rect 18550 23280 18590 23320
rect 18630 23280 18670 23320
rect 18710 23280 18750 23320
rect 18790 23280 18830 23320
rect 18870 23280 18910 23320
rect 18950 23280 18990 23320
rect 19030 23280 19070 23320
rect 19110 23280 19150 23320
rect 19190 23280 19230 23320
rect 19270 23280 19310 23320
rect 19350 23280 19390 23320
rect 19430 23280 19470 23320
rect 19510 23280 19550 23320
rect 19590 23280 19630 23320
rect 19670 23280 19710 23320
rect 19750 23280 19790 23320
rect 19830 23280 19870 23320
rect 19910 23280 19950 23320
rect 19990 23280 20030 23320
rect 20070 23280 20110 23320
rect 20150 23280 20190 23320
rect 20230 23280 20270 23320
rect 20310 23280 20350 23320
rect 20390 23280 20430 23320
rect 20470 23280 20510 23320
rect 20550 23280 20590 23320
rect 7640 22730 7680 22770
rect 7380 22640 7420 22680
rect 8650 22710 8690 22750
rect 9090 23080 9160 23140
rect 9100 22860 9150 22910
rect 9840 22730 9880 22770
rect 7880 22630 7920 22670
rect 7960 22630 8000 22670
rect 8260 22630 8300 22670
rect 8500 22630 8540 22670
rect 7480 22520 7520 22560
rect 7480 21660 7520 21700
rect 7740 22520 7780 22560
rect 7740 21640 7780 21680
rect 8800 22630 8840 22670
rect 8880 22630 8920 22670
rect 9000 22630 9040 22670
rect 9220 22640 9280 22700
rect 10410 22720 10480 22780
rect 10830 22730 10870 22770
rect 11410 22720 11480 22780
rect 11830 22730 11870 22770
rect 9580 22630 9620 22670
rect 10080 22620 10120 22660
rect 10160 22620 10200 22660
rect 10460 22620 10500 22660
rect 10570 22630 10610 22670
rect 11070 22620 11110 22660
rect 11150 22620 11190 22660
rect 11450 22620 11490 22660
rect 11570 22630 11610 22670
rect 12070 22620 12110 22660
rect 12150 22620 12190 22660
rect 12450 22620 12490 22660
rect 12530 22620 12570 22660
rect 12820 22630 12860 22670
rect 12900 22630 12940 22670
rect 13000 22630 13040 22670
rect 9680 22510 9720 22550
rect 9680 21630 9720 21670
rect 9940 22510 9980 22550
rect 9940 21630 9980 21670
rect 10670 22510 10710 22550
rect 10670 21630 10710 21670
rect 10930 22510 10970 22550
rect 10930 21630 10970 21670
rect 11670 22510 11710 22550
rect 11670 21630 11710 21670
rect 11930 22510 11970 22550
rect 11930 21630 11970 21670
rect 13130 22630 13170 22670
rect 13340 22630 13380 22670
rect 13230 22530 13270 22570
rect 13230 21640 13270 21680
rect 13470 22630 13510 22670
rect 13900 22630 13940 22670
rect 13570 22530 13610 22570
rect 13790 22530 13830 22570
rect 13570 21640 13610 21680
rect 13790 21640 13830 21680
rect 14030 22630 14070 22670
rect 14900 22630 14940 22670
rect 14130 22510 14170 22550
rect 14350 22510 14390 22550
rect 14570 22510 14610 22550
rect 14790 22510 14830 22550
rect 14130 21620 14170 21660
rect 14350 21620 14390 21660
rect 14570 21620 14610 21660
rect 14790 21620 14830 21660
rect 15090 22630 15130 22670
rect 16890 22630 16940 22680
rect 17040 22630 17080 22670
rect 15190 22510 15230 22550
rect 15410 22510 15450 22550
rect 15630 22510 15670 22550
rect 15850 22510 15890 22550
rect 16070 22510 16110 22550
rect 16290 22510 16330 22550
rect 16510 22510 16550 22550
rect 16730 22510 16770 22550
rect 15190 21620 15230 21660
rect 15410 21620 15450 21660
rect 15630 21620 15670 21660
rect 15850 21620 15890 21660
rect 16070 21620 16110 21660
rect 16290 21620 16330 21660
rect 16510 21620 16550 21660
rect 16730 21620 16770 21660
rect 20600 22630 20650 22680
rect 17140 22510 17180 22550
rect 17360 22510 17400 22550
rect 17580 22510 17620 22550
rect 17800 22510 17840 22550
rect 18020 22510 18060 22550
rect 18240 22510 18280 22550
rect 18460 22510 18500 22550
rect 18680 22510 18720 22550
rect 18900 22510 18940 22550
rect 19120 22510 19160 22550
rect 19340 22510 19380 22550
rect 19560 22510 19600 22550
rect 19780 22510 19820 22550
rect 20000 22510 20040 22550
rect 20220 22510 20260 22550
rect 20440 22510 20480 22550
rect 17140 21620 17180 21660
rect 17360 21620 17400 21660
rect 17580 21620 17620 21660
rect 17800 21620 17840 21660
rect 18020 21620 18060 21660
rect 18240 21620 18280 21660
rect 18460 21620 18500 21660
rect 18680 21620 18720 21660
rect 18900 21620 18940 21660
rect 19120 21620 19160 21660
rect 19340 21620 19380 21660
rect 19560 21620 19600 21660
rect 19780 21620 19820 21660
rect 20000 21620 20040 21660
rect 20220 21620 20260 21660
rect 20440 21620 20480 21660
rect 7320 20960 7360 21000
rect 7400 20960 7440 21000
rect 7480 20960 7520 21000
rect 7560 20960 7600 21000
rect 7640 20960 7680 21000
rect 7720 20960 7760 21000
rect 7800 20960 7840 21000
rect 7880 20960 7920 21000
rect 7960 20960 8000 21000
rect 8040 20960 8080 21000
rect 8120 20960 8160 21000
rect 8200 20960 8240 21000
rect 8280 20960 8320 21000
rect 8360 20960 8400 21000
rect 8440 20960 8480 21000
rect 8520 20960 8560 21000
rect 8600 20960 8640 21000
rect 8680 20960 8720 21000
rect 8760 20960 8800 21000
rect 8840 20960 8880 21000
rect 8920 20960 8960 21000
rect 9000 20960 9040 21000
rect 9080 20960 9120 21000
rect 9160 20960 9200 21000
rect 9260 20960 9300 21000
rect 9340 20960 9380 21000
rect 9420 20960 9460 21000
rect 9500 20960 9540 21000
rect 9580 20960 9620 21000
rect 9660 20960 9700 21000
rect 9740 20960 9780 21000
rect 9820 20960 9860 21000
rect 9900 20960 9940 21000
rect 9980 20960 10020 21000
rect 10060 20960 10100 21000
rect 10140 20960 10180 21000
rect 10220 20960 10260 21000
rect 10300 20960 10340 21000
rect 10380 20960 10420 21000
rect 10460 20960 10500 21000
rect 10540 20960 10580 21000
rect 10620 20960 10660 21000
rect 10700 20960 10740 21000
rect 10780 20960 10820 21000
rect 10860 20960 10900 21000
rect 10940 20960 10980 21000
rect 11020 20960 11060 21000
rect 11100 20960 11140 21000
rect 11180 20960 11220 21000
rect 11260 20960 11300 21000
rect 11340 20960 11380 21000
rect 11420 20960 11460 21000
rect 11500 20960 11540 21000
rect 11580 20960 11620 21000
rect 11660 20960 11700 21000
rect 11740 20960 11780 21000
rect 11820 20960 11860 21000
rect 11900 20960 11940 21000
rect 11980 20960 12020 21000
rect 12060 20960 12100 21000
rect 12140 20960 12180 21000
rect 12220 20960 12260 21000
rect 12300 20960 12340 21000
rect 12380 20960 12420 21000
rect 12460 20960 12500 21000
rect 12540 20960 12580 21000
rect 12620 20960 12660 21000
rect 12700 20960 12740 21000
rect 12780 20960 12820 21000
rect 12880 20960 12920 21000
rect 12960 20960 13000 21000
rect 13040 20960 13080 21000
rect 13120 20960 13160 21000
rect 13200 20960 13240 21000
rect 13280 20960 13320 21000
rect 13360 20960 13400 21000
rect 13440 20960 13480 21000
rect 13520 20960 13560 21000
rect 13600 20960 13640 21000
rect 13680 20960 13720 21000
rect 13760 20960 13800 21000
rect 13840 20960 13880 21000
rect 13920 20960 13960 21000
rect 14000 20960 14040 21000
rect 14080 20960 14120 21000
rect 14160 20960 14200 21000
rect 14240 20960 14280 21000
rect 14320 20960 14360 21000
rect 14400 20960 14440 21000
rect 14480 20960 14520 21000
rect 14560 20960 14600 21000
rect 14640 20960 14680 21000
rect 14720 20960 14760 21000
rect 14800 20960 14840 21000
rect 14880 20960 14920 21000
rect 14960 20960 15000 21000
rect 15040 20960 15080 21000
rect 15120 20960 15160 21000
rect 15200 20960 15240 21000
rect 15280 20960 15320 21000
rect 15360 20960 15400 21000
rect 15440 20960 15480 21000
rect 15520 20960 15560 21000
rect 15600 20960 15640 21000
rect 15680 20960 15720 21000
rect 15760 20960 15800 21000
rect 15840 20960 15880 21000
rect 15920 20960 15960 21000
rect 16000 20960 16040 21000
rect 16080 20960 16120 21000
rect 16160 20960 16200 21000
rect 16240 20960 16280 21000
rect 16320 20960 16360 21000
rect 16400 20960 16440 21000
rect 16480 20960 16520 21000
rect 16560 20960 16600 21000
rect 16640 20960 16680 21000
rect 16720 20960 16760 21000
rect 16800 20960 16840 21000
rect 16880 20960 16920 21000
rect 16960 20960 17000 21000
rect 17040 20960 17080 21000
rect 17120 20960 17160 21000
rect 17200 20960 17240 21000
rect 17280 20960 17320 21000
rect 17360 20960 17400 21000
rect 17440 20960 17480 21000
rect 17520 20960 17560 21000
rect 17600 20960 17640 21000
rect 17680 20960 17720 21000
rect 17760 20960 17800 21000
rect 17840 20960 17880 21000
rect 17920 20960 17960 21000
rect 18000 20960 18040 21000
rect 18080 20960 18120 21000
rect 18160 20960 18200 21000
rect 18240 20960 18280 21000
rect 18320 20960 18360 21000
rect 18400 20960 18440 21000
rect 18480 20960 18520 21000
rect 18560 20960 18600 21000
rect 18640 20960 18680 21000
rect 18720 20960 18760 21000
rect 18800 20960 18840 21000
rect 18880 20960 18920 21000
rect 18960 20960 19000 21000
rect 19040 20960 19080 21000
rect 19120 20960 19160 21000
rect 19200 20960 19240 21000
rect 19280 20960 19320 21000
rect 19360 20960 19400 21000
rect 19440 20960 19480 21000
rect 19520 20960 19560 21000
rect 19600 20960 19640 21000
rect 19680 20960 19720 21000
rect 19760 20960 19800 21000
rect 19840 20960 19880 21000
rect 19920 20960 19960 21000
rect 20000 20960 20040 21000
rect 20080 20960 20120 21000
rect 20160 20960 20200 21000
rect 20240 20960 20280 21000
rect 20320 20960 20360 21000
rect 20400 20960 20440 21000
rect 20480 20960 20520 21000
rect 20560 20960 20600 21000
rect 7320 20430 7360 20470
rect 7400 20430 7440 20470
rect 7480 20430 7520 20470
rect 7560 20430 7600 20470
rect 7640 20430 7680 20470
rect 7720 20430 7760 20470
rect 7800 20430 7840 20470
rect 7880 20430 7920 20470
rect 7960 20430 8000 20470
rect 8040 20430 8080 20470
rect 8120 20430 8160 20470
rect 7110 19410 7170 19470
rect 7400 19270 7440 19310
rect 6960 18620 7020 18680
rect 7230 18360 7290 18420
rect 7400 18390 7440 18430
rect 12730 20350 12800 20410
rect 8360 19980 8400 20020
rect 8440 19980 8480 20020
rect 8520 19980 8560 20020
rect 8600 19980 8640 20020
rect 8680 19980 8720 20020
rect 8760 19980 8800 20020
rect 8840 19980 8880 20020
rect 8920 19980 8960 20020
rect 9000 19980 9040 20020
rect 9080 19980 9120 20020
rect 9160 19980 9200 20020
rect 9260 19980 9300 20020
rect 9340 19980 9380 20020
rect 9420 19980 9460 20020
rect 9500 19980 9540 20020
rect 9580 19980 9620 20020
rect 9660 19980 9700 20020
rect 9740 19980 9780 20020
rect 9820 19980 9860 20020
rect 9900 19980 9940 20020
rect 9980 19980 10020 20020
rect 10060 19980 10100 20020
rect 10140 19980 10180 20020
rect 10220 19980 10260 20020
rect 10300 19980 10340 20020
rect 10380 19980 10420 20020
rect 10460 19980 10500 20020
rect 10540 19980 10580 20020
rect 10620 19980 10660 20020
rect 10700 19980 10740 20020
rect 10780 19980 10820 20020
rect 10860 19980 10900 20020
rect 10940 19980 10980 20020
rect 11020 19980 11060 20020
rect 11100 19980 11140 20020
rect 11180 19980 11220 20020
rect 11260 19980 11300 20020
rect 11340 19980 11380 20020
rect 11420 19980 11460 20020
rect 11500 19980 11540 20020
rect 11580 19980 11620 20020
rect 11660 19980 11700 20020
rect 11740 19980 11780 20020
rect 11820 19980 11860 20020
rect 11900 19980 11940 20020
rect 11980 19980 12020 20020
rect 12060 19980 12100 20020
rect 12140 19980 12180 20020
rect 12220 19980 12260 20020
rect 12300 19980 12340 20020
rect 12380 19980 12420 20020
rect 12460 19980 12500 20020
rect 12540 19980 12580 20020
rect 12620 19980 12660 20020
rect 12700 19980 12740 20020
rect 12780 19980 12820 20020
rect 12860 19980 12900 20020
rect 12940 19980 12980 20020
rect 13040 19980 13080 20020
rect 13120 19980 13160 20020
rect 13200 19980 13240 20020
rect 13280 19980 13320 20020
rect 13360 19980 13400 20020
rect 13440 19980 13480 20020
rect 13520 19980 13560 20020
rect 13600 19980 13640 20020
rect 13680 19980 13720 20020
rect 13760 19980 13800 20020
rect 13840 19980 13880 20020
rect 13920 19980 13960 20020
rect 14000 19980 14040 20020
rect 14080 19980 14120 20020
rect 14160 19980 14200 20020
rect 14240 19980 14280 20020
rect 14320 19980 14360 20020
rect 14400 19980 14440 20020
rect 14480 19980 14520 20020
rect 14560 19980 14600 20020
rect 14640 19980 14680 20020
rect 14720 19980 14760 20020
rect 14800 19980 14840 20020
rect 14880 19980 14920 20020
rect 14960 19980 15000 20020
rect 15040 19980 15080 20020
rect 15120 19980 15160 20020
rect 15200 19980 15240 20020
rect 15280 19980 15320 20020
rect 15360 19980 15400 20020
rect 15440 19980 15480 20020
rect 15520 19980 15560 20020
rect 15600 19980 15640 20020
rect 15680 19980 15720 20020
rect 15760 19980 15800 20020
rect 15840 19980 15880 20020
rect 15920 19980 15960 20020
rect 16000 19980 16040 20020
rect 16080 19980 16120 20020
rect 16160 19980 16200 20020
rect 16240 19980 16280 20020
rect 16320 19980 16360 20020
rect 16400 19980 16440 20020
rect 16480 19980 16520 20020
rect 16560 19980 16600 20020
rect 16640 19980 16680 20020
rect 16720 19980 16760 20020
rect 16800 19980 16840 20020
rect 16880 19980 16920 20020
rect 16960 19980 17000 20020
rect 17040 19980 17080 20020
rect 17120 19980 17160 20020
rect 17200 19980 17240 20020
rect 17280 19980 17320 20020
rect 17360 19980 17400 20020
rect 17440 19980 17480 20020
rect 17520 19980 17560 20020
rect 17600 19980 17640 20020
rect 17680 19980 17720 20020
rect 17760 19980 17800 20020
rect 17840 19980 17880 20020
rect 17920 19980 17960 20020
rect 18000 19980 18040 20020
rect 18080 19980 18120 20020
rect 18160 19980 18200 20020
rect 18240 19980 18280 20020
rect 18320 19980 18360 20020
rect 18400 19980 18440 20020
rect 18480 19980 18520 20020
rect 18560 19980 18600 20020
rect 18640 19980 18680 20020
rect 18720 19980 18760 20020
rect 18800 19980 18840 20020
rect 18880 19980 18920 20020
rect 18960 19980 19000 20020
rect 19040 19980 19080 20020
rect 19120 19980 19160 20020
rect 19200 19980 19240 20020
rect 19280 19980 19320 20020
rect 19360 19980 19400 20020
rect 19440 19980 19480 20020
rect 19520 19980 19560 20020
rect 19600 19980 19640 20020
rect 19680 19980 19720 20020
rect 19760 19980 19800 20020
rect 19840 19980 19880 20020
rect 19920 19980 19960 20020
rect 20000 19980 20040 20020
rect 20080 19980 20120 20020
rect 20160 19980 20200 20020
rect 20240 19980 20280 20020
rect 20320 19980 20360 20020
rect 20400 19980 20440 20020
rect 20480 19980 20520 20020
rect 20560 19980 20600 20020
rect 7560 18240 7600 18280
rect 7300 18130 7340 18170
rect 7970 18240 8010 18280
rect 8500 18310 8540 18350
rect 8800 18310 8840 18350
rect 8880 18310 8920 18350
rect 9000 18310 9040 18350
rect 8650 18230 8690 18270
rect 7780 18030 7820 18070
rect 8190 18030 8230 18070
rect 9220 18270 9280 18330
rect 9680 19320 9720 19360
rect 9680 18430 9720 18470
rect 9940 19320 9980 19360
rect 9940 18430 9980 18470
rect 10670 19320 10710 19360
rect 10670 18430 10710 18470
rect 10930 19320 10970 19360
rect 10930 18430 10970 18470
rect 11670 19310 11710 19350
rect 11670 18420 11710 18460
rect 11930 19310 11970 19350
rect 11930 18420 11970 18460
rect 9580 18310 9620 18350
rect 10080 18320 10120 18360
rect 10160 18320 10200 18360
rect 10460 18320 10500 18360
rect 10570 18310 10610 18350
rect 11070 18320 11110 18360
rect 11150 18320 11190 18360
rect 11450 18320 11490 18360
rect 11570 18310 11610 18350
rect 12070 18320 12110 18360
rect 12150 18320 12190 18360
rect 12450 18320 12490 18360
rect 12530 18320 12570 18360
rect 12820 18310 12860 18350
rect 12900 18310 12940 18350
rect 9840 18210 9880 18250
rect 9100 18130 9150 18180
rect 9090 17900 9160 17960
rect 9470 18040 9540 18100
rect 10410 18200 10480 18260
rect 10830 18210 10870 18250
rect 11830 18210 11870 18250
rect 13230 19300 13270 19340
rect 13230 18410 13270 18450
rect 13000 18310 13040 18350
rect 13130 18310 13170 18350
rect 13570 19300 13610 19340
rect 13790 19300 13830 19340
rect 13570 18410 13610 18450
rect 13790 18410 13830 18450
rect 13340 18310 13380 18350
rect 13470 18310 13510 18350
rect 14130 19320 14170 19360
rect 14350 19320 14390 19360
rect 14570 19320 14610 19360
rect 14790 19320 14830 19360
rect 14130 18430 14170 18470
rect 14350 18430 14390 18470
rect 14570 18430 14610 18470
rect 14790 18430 14830 18470
rect 13900 18310 13940 18350
rect 14030 18310 14070 18350
rect 15190 19320 15230 19360
rect 15410 19320 15450 19360
rect 15630 19320 15670 19360
rect 15850 19320 15890 19360
rect 16070 19320 16110 19360
rect 16290 19320 16330 19360
rect 16510 19320 16550 19360
rect 16730 19320 16770 19360
rect 15190 18430 15230 18470
rect 15410 18430 15450 18470
rect 15630 18430 15670 18470
rect 15850 18430 15890 18470
rect 16070 18430 16110 18470
rect 16290 18430 16330 18470
rect 16510 18430 16550 18470
rect 16730 18430 16770 18470
rect 14900 18310 14940 18350
rect 15090 18310 15130 18350
rect 17140 19320 17180 19360
rect 17360 19320 17400 19360
rect 17580 19320 17620 19360
rect 17800 19320 17840 19360
rect 18020 19320 18060 19360
rect 18240 19320 18280 19360
rect 18460 19320 18500 19360
rect 18680 19320 18720 19360
rect 18900 19320 18940 19360
rect 19120 19320 19160 19360
rect 19340 19320 19380 19360
rect 19560 19320 19600 19360
rect 19780 19320 19820 19360
rect 20000 19320 20040 19360
rect 20220 19320 20260 19360
rect 20440 19320 20480 19360
rect 17140 18430 17180 18470
rect 17360 18430 17400 18470
rect 17580 18430 17620 18470
rect 17800 18430 17840 18470
rect 18020 18430 18060 18470
rect 18240 18430 18280 18470
rect 18460 18430 18500 18470
rect 18680 18430 18720 18470
rect 18900 18430 18940 18470
rect 19120 18430 19160 18470
rect 19340 18430 19380 18470
rect 19560 18430 19600 18470
rect 19780 18430 19820 18470
rect 20000 18430 20040 18470
rect 20220 18430 20260 18470
rect 20440 18430 20480 18470
rect 16890 18300 16940 18350
rect 17040 18310 17080 18350
rect 20600 18300 20650 18350
rect 7320 17660 7360 17700
rect 7400 17660 7440 17700
rect 7480 17660 7520 17700
rect 7560 17660 7600 17700
rect 7640 17660 7680 17700
rect 7720 17660 7760 17700
rect 7800 17660 7840 17700
rect 7880 17660 7920 17700
rect 7960 17660 8000 17700
rect 8040 17660 8080 17700
rect 8120 17660 8160 17700
rect 8200 17660 8240 17700
rect 8280 17660 8320 17700
rect 8360 17660 8400 17700
rect 8440 17660 8480 17700
rect 8520 17660 8560 17700
rect 8600 17660 8640 17700
rect 8680 17660 8720 17700
rect 8760 17660 8800 17700
rect 8840 17660 8880 17700
rect 8920 17660 8960 17700
rect 9000 17660 9040 17700
rect 9080 17660 9120 17700
rect 9160 17660 9200 17700
rect 9270 17660 9310 17700
rect 9350 17660 9390 17700
rect 9430 17660 9470 17700
rect 9510 17660 9550 17700
rect 9590 17660 9630 17700
rect 9670 17660 9710 17700
rect 9750 17660 9790 17700
rect 9830 17660 9870 17700
rect 9910 17660 9950 17700
rect 9990 17660 10030 17700
rect 10070 17660 10110 17700
rect 10150 17660 10190 17700
rect 10230 17660 10270 17700
rect 10310 17660 10350 17700
rect 10390 17660 10430 17700
rect 10470 17660 10510 17700
rect 10550 17660 10590 17700
rect 10630 17660 10670 17700
rect 10710 17660 10750 17700
rect 10790 17660 10830 17700
rect 10870 17660 10910 17700
rect 10950 17660 10990 17700
rect 11030 17660 11070 17700
rect 11110 17660 11150 17700
rect 11190 17660 11230 17700
rect 11270 17660 11310 17700
rect 11350 17660 11390 17700
rect 11430 17660 11470 17700
rect 11510 17660 11550 17700
rect 11590 17660 11630 17700
rect 11670 17660 11710 17700
rect 11750 17660 11790 17700
rect 11830 17660 11870 17700
rect 11910 17660 11950 17700
rect 11990 17660 12030 17700
rect 12070 17660 12110 17700
rect 12150 17660 12190 17700
rect 12230 17660 12270 17700
rect 12310 17660 12350 17700
rect 12390 17660 12430 17700
rect 12470 17660 12510 17700
rect 12550 17660 12590 17700
rect 12630 17660 12670 17700
rect 12710 17660 12750 17700
rect 12790 17660 12830 17700
rect 12870 17660 12910 17700
rect 12950 17660 12990 17700
rect 13030 17660 13070 17700
rect 13110 17660 13150 17700
rect 13190 17660 13230 17700
rect 13270 17660 13310 17700
rect 13350 17660 13390 17700
rect 13430 17660 13470 17700
rect 13510 17660 13550 17700
rect 13590 17660 13630 17700
rect 13670 17660 13710 17700
rect 13750 17660 13790 17700
rect 13830 17660 13870 17700
rect 13910 17660 13950 17700
rect 13990 17660 14030 17700
rect 14070 17660 14110 17700
rect 14150 17660 14190 17700
rect 14230 17660 14270 17700
rect 14310 17660 14350 17700
rect 14390 17660 14430 17700
rect 14470 17660 14510 17700
rect 14550 17660 14590 17700
rect 14630 17660 14670 17700
rect 14710 17660 14750 17700
rect 14790 17660 14830 17700
rect 14870 17660 14910 17700
rect 14950 17660 14990 17700
rect 15030 17660 15070 17700
rect 15110 17660 15150 17700
rect 15190 17660 15230 17700
rect 15270 17660 15310 17700
rect 15350 17660 15390 17700
rect 15430 17660 15470 17700
rect 15510 17660 15550 17700
rect 15590 17660 15630 17700
rect 15670 17660 15710 17700
rect 15750 17660 15790 17700
rect 15830 17660 15870 17700
rect 15910 17660 15950 17700
rect 15990 17660 16030 17700
rect 16070 17660 16110 17700
rect 16150 17660 16190 17700
rect 16230 17660 16270 17700
rect 16310 17660 16350 17700
rect 16390 17660 16430 17700
rect 16470 17660 16510 17700
rect 16550 17660 16590 17700
rect 16630 17660 16670 17700
rect 16710 17660 16750 17700
rect 16790 17660 16830 17700
rect 16870 17660 16910 17700
rect 16950 17660 16990 17700
rect 17030 17660 17070 17700
rect 17110 17660 17150 17700
rect 17190 17660 17230 17700
rect 17270 17660 17310 17700
rect 17350 17660 17390 17700
rect 17430 17660 17470 17700
rect 17510 17660 17550 17700
rect 17590 17660 17630 17700
rect 17670 17660 17710 17700
rect 17750 17660 17790 17700
rect 17830 17660 17870 17700
rect 17910 17660 17950 17700
rect 17990 17660 18030 17700
rect 18070 17660 18110 17700
rect 18150 17660 18190 17700
rect 18230 17660 18270 17700
rect 18310 17660 18350 17700
rect 18390 17660 18430 17700
rect 18470 17660 18510 17700
rect 18550 17660 18590 17700
rect 18630 17660 18670 17700
rect 18710 17660 18750 17700
rect 18790 17660 18830 17700
rect 18870 17660 18910 17700
rect 18950 17660 18990 17700
rect 19030 17660 19070 17700
rect 19110 17660 19150 17700
rect 19190 17660 19230 17700
rect 19270 17660 19310 17700
rect 19350 17660 19390 17700
rect 19430 17660 19470 17700
rect 19510 17660 19550 17700
rect 19590 17660 19630 17700
rect 19670 17660 19710 17700
rect 19750 17660 19790 17700
rect 19830 17660 19870 17700
rect 19910 17660 19950 17700
rect 19990 17660 20030 17700
rect 20070 17660 20110 17700
rect 20150 17660 20190 17700
rect 20230 17660 20270 17700
rect 20310 17660 20350 17700
rect 20390 17660 20430 17700
rect 20470 17660 20510 17700
rect 20550 17660 20590 17700
rect 9710 15620 9750 15660
rect 9790 15620 9830 15660
rect 9870 15620 9910 15660
rect 9950 15620 9990 15660
rect 10030 15620 10070 15660
rect 10110 15620 10150 15660
rect 10190 15620 10230 15660
rect 10270 15620 10310 15660
rect 10350 15620 10390 15660
rect 10430 15620 10470 15660
rect 10510 15620 10550 15660
rect 10590 15620 10630 15660
rect 10670 15620 10710 15660
rect 10750 15620 10790 15660
rect 10830 15620 10870 15660
rect 10910 15620 10950 15660
rect 10990 15620 11030 15660
rect 11070 15620 11110 15660
rect 11150 15620 11190 15660
rect 11230 15620 11270 15660
rect 11310 15620 11350 15660
rect 11390 15620 11430 15660
rect 11470 15620 11510 15660
rect 11550 15620 11590 15660
rect 11630 15620 11670 15660
rect 11710 15620 11750 15660
rect 11790 15620 11830 15660
rect 11870 15620 11910 15660
rect 11950 15620 11990 15660
rect 12030 15620 12070 15660
rect 12110 15620 12150 15660
rect 12190 15620 12230 15660
rect 12270 15620 12310 15660
rect 12350 15620 12390 15660
rect 12430 15620 12470 15660
rect 12510 15620 12550 15660
rect 12590 15620 12630 15660
rect 12670 15620 12710 15660
rect 12750 15620 12790 15660
rect 12830 15620 12870 15660
rect 12910 15620 12950 15660
rect 12990 15620 13030 15660
rect 13070 15620 13110 15660
rect 13150 15620 13190 15660
rect 13230 15620 13270 15660
rect 13310 15620 13350 15660
rect 13390 15620 13430 15660
rect 13470 15620 13510 15660
rect 13550 15620 13590 15660
rect 13630 15620 13670 15660
rect 13710 15620 13750 15660
rect 13790 15620 13830 15660
rect 13870 15620 13910 15660
rect 13950 15620 13990 15660
rect 14030 15620 14070 15660
rect 14110 15620 14150 15660
rect 14190 15620 14230 15660
rect 14270 15620 14310 15660
rect 14350 15620 14390 15660
rect 14430 15620 14470 15660
rect 14510 15620 14550 15660
rect 14590 15620 14630 15660
rect 14670 15620 14710 15660
rect 14750 15620 14790 15660
rect 14830 15620 14870 15660
rect 14910 15620 14950 15660
rect 14990 15620 15030 15660
rect 15070 15620 15110 15660
rect 15150 15620 15190 15660
rect 15230 15620 15270 15660
rect 15310 15620 15350 15660
rect 15390 15620 15430 15660
rect 15470 15620 15510 15660
rect 15550 15620 15590 15660
rect 15630 15620 15670 15660
rect 15710 15620 15750 15660
rect 15790 15620 15830 15660
rect 15870 15620 15910 15660
rect 15950 15620 15990 15660
rect 16030 15620 16070 15660
rect 16110 15620 16150 15660
rect 16190 15620 16230 15660
rect 16270 15620 16310 15660
rect 16350 15620 16390 15660
rect 16430 15620 16470 15660
rect 16510 15620 16550 15660
rect 16590 15620 16630 15660
rect 16670 15620 16710 15660
rect 16750 15620 16790 15660
rect 16830 15620 16870 15660
rect 16910 15620 16950 15660
rect 16990 15620 17030 15660
rect 17070 15620 17110 15660
rect 17150 15620 17190 15660
rect 17230 15620 17270 15660
rect 17310 15620 17350 15660
rect 17390 15620 17430 15660
rect 17470 15620 17510 15660
rect 17550 15620 17590 15660
rect 17630 15620 17670 15660
rect 17710 15620 17750 15660
rect 17790 15620 17830 15660
rect 17870 15620 17910 15660
rect 17950 15620 17990 15660
rect 18030 15620 18070 15660
rect 18110 15620 18150 15660
rect 18190 15620 18230 15660
rect 18270 15620 18310 15660
rect 18350 15620 18390 15660
rect 18430 15620 18470 15660
rect 18510 15620 18550 15660
rect 18590 15620 18630 15660
rect 18670 15620 18710 15660
rect 18750 15620 18790 15660
rect 18830 15620 18870 15660
rect 18910 15620 18950 15660
rect 18990 15620 19030 15660
rect 19070 15620 19110 15660
rect 19150 15620 19190 15660
rect 19230 15620 19270 15660
rect 19310 15620 19350 15660
rect 19390 15620 19430 15660
rect 19470 15620 19510 15660
rect 19550 15620 19590 15660
rect 19630 15620 19670 15660
rect 19710 15620 19750 15660
rect 19800 15620 19840 15660
rect 19880 15620 19920 15660
rect 19960 15620 20000 15660
rect 20040 15620 20080 15660
rect 20120 15620 20160 15660
rect 20200 15620 20240 15660
rect 20280 15620 20320 15660
rect 20370 15620 20410 15660
rect 20450 15620 20490 15660
rect 20530 15620 20570 15660
rect 20610 15620 20650 15660
rect 20690 15620 20730 15660
rect 20770 15620 20810 15660
rect 20850 15620 20890 15660
rect 20930 15620 20970 15660
rect 21010 15620 21050 15660
rect 21090 15620 21130 15660
rect 7430 15230 7500 15290
rect 9750 15050 9810 15110
rect 10580 15070 10620 15110
rect 10060 14960 10100 15000
rect 10280 14960 10350 15020
rect 11570 15070 11610 15110
rect 12570 15070 12610 15110
rect 10820 14960 10860 15000
rect 10900 14960 10940 15000
rect 11200 14960 11240 15000
rect 11310 14970 11350 15010
rect 11810 14960 11850 15000
rect 11890 14960 11930 15000
rect 12190 14960 12230 15000
rect 12310 14970 12350 15010
rect 12810 14960 12850 15000
rect 12890 14960 12930 15000
rect 13180 14970 13220 15010
rect 13260 14970 13300 15010
rect 13360 14970 13400 15010
rect 13490 14970 13530 15010
rect 13700 14970 13740 15010
rect 13830 14970 13870 15010
rect 14260 14970 14300 15010
rect 14390 14970 14430 15010
rect 15260 14970 15300 15010
rect 15450 14970 15490 15010
rect 17250 14970 17300 15020
rect 17400 14970 17440 15010
rect 20960 14970 21010 15020
rect 9700 14300 9740 14340
rect 9790 14300 9830 14340
rect 9870 14300 9910 14340
rect 9950 14300 9990 14340
rect 10030 14300 10070 14340
rect 10110 14300 10150 14340
rect 10190 14300 10230 14340
rect 10270 14300 10310 14340
rect 10350 14300 10390 14340
rect 10430 14300 10470 14340
rect 10510 14300 10550 14340
rect 10590 14300 10630 14340
rect 10670 14300 10710 14340
rect 10750 14300 10790 14340
rect 10830 14300 10870 14340
rect 10910 14300 10950 14340
rect 10990 14300 11030 14340
rect 11070 14300 11110 14340
rect 11150 14300 11190 14340
rect 11230 14300 11270 14340
rect 11310 14300 11350 14340
rect 11390 14300 11430 14340
rect 11470 14300 11510 14340
rect 11550 14300 11590 14340
rect 11630 14300 11670 14340
rect 11710 14300 11750 14340
rect 11790 14300 11830 14340
rect 11870 14300 11910 14340
rect 11950 14300 11990 14340
rect 12030 14300 12070 14340
rect 12110 14300 12150 14340
rect 12190 14300 12230 14340
rect 12270 14300 12310 14340
rect 12350 14300 12390 14340
rect 12430 14300 12470 14340
rect 12510 14300 12550 14340
rect 12590 14300 12630 14340
rect 12670 14300 12710 14340
rect 12750 14300 12790 14340
rect 12830 14300 12870 14340
rect 12910 14300 12950 14340
rect 12990 14300 13030 14340
rect 13070 14300 13110 14340
rect 13150 14300 13230 14340
rect 13270 14300 13310 14340
rect 13350 14300 13390 14340
rect 13430 14300 13470 14340
rect 13510 14300 13550 14340
rect 13590 14300 13630 14340
rect 13670 14300 13710 14340
rect 13750 14300 13790 14340
rect 13830 14300 13870 14340
rect 13910 14300 13950 14340
rect 13990 14300 14030 14340
rect 14070 14300 14110 14340
rect 14150 14300 14190 14340
rect 14230 14300 14270 14340
rect 14310 14300 14350 14340
rect 14390 14300 14430 14340
rect 14470 14300 14510 14340
rect 14550 14300 14590 14340
rect 14630 14300 14670 14340
rect 14710 14300 14750 14340
rect 14790 14300 14830 14340
rect 14870 14300 14910 14340
rect 14950 14300 14990 14340
rect 15030 14300 15070 14340
rect 15110 14300 15150 14340
rect 15190 14300 15230 14340
rect 15270 14300 15310 14340
rect 15350 14300 15390 14340
rect 15430 14300 15470 14340
rect 15510 14300 15550 14340
rect 15590 14300 15630 14340
rect 15670 14300 15710 14340
rect 15750 14300 15790 14340
rect 15830 14300 15870 14340
rect 15910 14300 15950 14340
rect 15990 14300 16030 14340
rect 16070 14300 16110 14340
rect 16150 14300 16190 14340
rect 16230 14300 16270 14340
rect 16310 14300 16350 14340
rect 16390 14300 16430 14340
rect 16470 14300 16510 14340
rect 16550 14300 16590 14340
rect 16630 14300 16670 14340
rect 16710 14300 16750 14340
rect 16790 14300 16830 14340
rect 16870 14300 16910 14340
rect 16950 14300 16990 14340
rect 17030 14300 17070 14340
rect 17110 14300 17150 14340
rect 17190 14300 17230 14340
rect 17270 14300 17310 14340
rect 17350 14300 17390 14340
rect 17430 14300 17470 14340
rect 17510 14300 17550 14340
rect 17590 14300 17630 14340
rect 17670 14300 17710 14340
rect 17750 14300 17790 14340
rect 17830 14300 17870 14340
rect 17910 14300 17950 14340
rect 17990 14300 18030 14340
rect 18070 14300 18110 14340
rect 18150 14300 18190 14340
rect 18230 14300 18270 14340
rect 18310 14300 18350 14340
rect 18390 14300 18430 14340
rect 18470 14300 18510 14340
rect 18550 14300 18590 14340
rect 18630 14300 18670 14340
rect 18710 14300 18750 14340
rect 18790 14300 18830 14340
rect 18870 14300 18910 14340
rect 18950 14300 18990 14340
rect 19030 14300 19070 14340
rect 19110 14300 19150 14340
rect 19190 14300 19230 14340
rect 19270 14300 19310 14340
rect 19350 14300 19390 14340
rect 19430 14300 19470 14340
rect 19510 14300 19550 14340
rect 19590 14300 19630 14340
rect 19670 14300 19710 14340
rect 19750 14300 19790 14340
rect 19830 14300 19870 14340
rect 19910 14300 19950 14340
rect 19990 14300 20030 14340
rect 20070 14300 20110 14340
rect 20150 14300 20190 14340
rect 20230 14300 20270 14340
rect 20310 14300 20350 14340
rect 20390 14300 20430 14340
rect 20470 14300 20510 14340
rect 20550 14300 20590 14340
rect 20630 14300 20670 14340
rect 20710 14300 20750 14340
rect 20790 14300 20830 14340
rect 20870 14300 20910 14340
rect 20950 14300 20990 14340
rect 21030 14300 21070 14340
rect 8430 14200 8500 14260
rect 7320 13330 7360 13370
rect 7400 13330 7440 13370
rect 7480 13330 7520 13370
rect 7560 13330 7600 13370
rect 7640 13330 7680 13370
rect 7720 13330 7760 13370
rect 7800 13330 7840 13370
rect 7880 13330 7920 13370
rect 7960 13330 8000 13370
rect 8040 13330 8080 13370
rect 8120 13330 8160 13370
rect 8200 13330 8240 13370
rect 8280 13330 8320 13370
rect 8360 13330 8400 13370
rect 8440 13330 8480 13370
rect 8520 13330 8560 13370
rect 8600 13330 8640 13370
rect 8680 13330 8720 13370
rect 8760 13330 8800 13370
rect 8840 13330 8880 13370
rect 8920 13330 8960 13370
rect 9000 13330 9040 13370
rect 9080 13330 9120 13370
rect 9160 13330 9200 13370
rect 9240 13330 9280 13370
rect 9320 13330 9360 13370
rect 9400 13330 9440 13370
rect 9480 13330 9520 13370
rect 9560 13330 9600 13370
rect 9640 13330 9680 13370
rect 9720 13330 9760 13370
rect 9800 13330 9840 13370
rect 9890 13330 9930 13370
rect 9970 13330 10010 13370
rect 10050 13330 10090 13370
rect 10130 13330 10170 13370
rect 10210 13330 10250 13370
rect 10290 13330 10330 13370
rect 10370 13330 10410 13370
rect 10450 13330 10490 13370
rect 10530 13330 10570 13370
rect 10610 13330 10650 13370
rect 10690 13330 10730 13370
rect 10770 13330 10810 13370
rect 10850 13330 10890 13370
rect 10930 13330 10970 13370
rect 11010 13330 11050 13370
rect 11090 13330 11130 13370
rect 11170 13330 11210 13370
rect 11250 13330 11290 13370
rect 11330 13330 11370 13370
rect 11410 13330 11450 13370
rect 11490 13330 11530 13370
rect 11570 13330 11610 13370
rect 11650 13330 11690 13370
rect 11730 13330 11770 13370
rect 11810 13330 11850 13370
rect 11890 13330 11930 13370
rect 11970 13330 12010 13370
rect 12050 13330 12090 13370
rect 12130 13330 12170 13370
rect 12210 13330 12250 13370
rect 12290 13330 12330 13370
rect 12370 13330 12410 13370
rect 12450 13330 12490 13370
rect 12530 13330 12570 13370
rect 12610 13330 12650 13370
rect 12690 13330 12730 13370
rect 12770 13330 12810 13370
rect 12850 13330 12890 13370
rect 12930 13330 12970 13370
rect 13010 13330 13050 13370
rect 13090 13330 13130 13370
rect 13170 13330 13210 13370
rect 13250 13330 13290 13370
rect 13330 13330 13400 13370
rect 13440 13330 13480 13370
rect 13520 13330 13560 13370
rect 13600 13330 13640 13370
rect 13680 13330 13720 13370
rect 13760 13330 13800 13370
rect 13840 13330 13880 13370
rect 13920 13330 13960 13370
rect 14000 13330 14040 13370
rect 14080 13330 14120 13370
rect 14160 13330 14200 13370
rect 14240 13330 14280 13370
rect 14320 13330 14360 13370
rect 14400 13330 14440 13370
rect 14480 13330 14520 13370
rect 14560 13330 14600 13370
rect 14640 13330 14680 13370
rect 14720 13330 14760 13370
rect 14800 13330 14840 13370
rect 14880 13330 14920 13370
rect 14960 13330 15000 13370
rect 15040 13330 15080 13370
rect 15120 13330 15160 13370
rect 15200 13330 15240 13370
rect 15280 13330 15320 13370
rect 15360 13330 15400 13370
rect 15440 13330 15480 13370
rect 15520 13330 15560 13370
rect 15600 13330 15640 13370
rect 15680 13330 15720 13370
rect 15760 13330 15800 13370
rect 15840 13330 15880 13370
rect 15920 13330 15960 13370
rect 16000 13330 16040 13370
rect 16080 13330 16120 13370
rect 16160 13330 16200 13370
rect 16240 13330 16280 13370
rect 16320 13330 16360 13370
rect 16400 13330 16440 13370
rect 16480 13330 16520 13370
rect 16560 13330 16600 13370
rect 16640 13330 16680 13370
rect 16720 13330 16760 13370
rect 16800 13330 16840 13370
rect 16880 13330 16920 13370
rect 16960 13330 17000 13370
rect 17040 13330 17080 13370
rect 17120 13330 17160 13370
rect 17200 13330 17240 13370
rect 17280 13330 17320 13370
rect 17360 13330 17400 13370
rect 17440 13330 17480 13370
rect 17520 13330 17560 13370
rect 17600 13330 17640 13370
rect 17680 13330 17720 13370
rect 17760 13330 17800 13370
rect 17840 13330 17880 13370
rect 17920 13330 17960 13370
rect 18000 13330 18040 13370
rect 18080 13330 18120 13370
rect 18160 13330 18200 13370
rect 18240 13330 18280 13370
rect 18320 13330 18360 13370
rect 18400 13330 18440 13370
rect 18480 13330 18520 13370
rect 18560 13330 18600 13370
rect 18640 13330 18680 13370
rect 18720 13330 18760 13370
rect 18800 13330 18840 13370
rect 18880 13330 18920 13370
rect 18960 13330 19000 13370
rect 19040 13330 19080 13370
rect 19120 13330 19160 13370
rect 19200 13330 19240 13370
rect 19280 13330 19320 13370
rect 19360 13330 19400 13370
rect 19440 13330 19480 13370
rect 19520 13330 19560 13370
rect 19600 13330 19640 13370
rect 19680 13330 19720 13370
rect 19760 13330 19800 13370
rect 19840 13330 19880 13370
rect 19920 13330 19960 13370
rect 20000 13330 20040 13370
rect 20080 13330 20120 13370
rect 20160 13330 20200 13370
rect 20240 13330 20280 13370
rect 20320 13330 20360 13370
rect 20400 13330 20440 13370
rect 20480 13330 20520 13370
rect 20560 13330 20600 13370
rect 20640 13330 20680 13370
rect 20720 13330 20760 13370
rect 20800 13330 20840 13370
rect 20880 13330 20920 13370
rect 20960 13330 21000 13370
rect 21040 13330 21080 13370
rect 9670 13090 9740 13150
rect 7270 12650 7330 12710
rect 7570 12660 7610 12700
rect 7700 12650 7760 12710
rect 7820 12660 7860 12700
rect 8320 12670 8360 12710
rect 7590 12540 7650 12600
rect 8080 12560 8120 12600
rect 8570 12650 8610 12690
rect 8870 12660 8910 12700
rect 8950 12660 8990 12700
rect 9070 12660 9110 12700
rect 9210 12660 9250 12700
rect 9330 12660 9370 12700
rect 9460 12660 9500 12700
rect 9580 12660 9620 12700
rect 9860 12670 9900 12710
rect 10160 12670 10200 12710
rect 10420 12660 10460 12700
rect 10920 12670 10960 12710
rect 11000 12670 11040 12710
rect 11300 12670 11340 12710
rect 11410 12660 11450 12700
rect 11910 12670 11950 12710
rect 11990 12670 12030 12710
rect 12290 12670 12330 12710
rect 12410 12660 12450 12700
rect 12910 12670 12950 12710
rect 12990 12670 13030 12710
rect 13280 12660 13320 12700
rect 13360 12660 13400 12700
rect 8720 12540 8760 12580
rect 9750 12470 9820 12530
rect 10680 12560 10720 12600
rect 11280 12550 11350 12610
rect 11670 12560 11710 12600
rect 12670 12560 12710 12600
rect 13460 12660 13500 12700
rect 13590 12660 13630 12700
rect 13800 12660 13840 12700
rect 13930 12660 13970 12700
rect 14360 12660 14400 12700
rect 14490 12660 14530 12700
rect 15360 12660 15400 12700
rect 15550 12660 15590 12700
rect 17350 12650 17400 12700
rect 17500 12660 17540 12700
rect 21060 12650 21110 12700
rect 9810 12010 9850 12050
rect 9890 12010 9930 12050
rect 9970 12010 10010 12050
rect 10050 12010 10090 12050
rect 10130 12010 10170 12050
rect 10210 12010 10250 12050
rect 10290 12010 10330 12050
rect 10370 12010 10410 12050
rect 10450 12010 10490 12050
rect 10530 12010 10570 12050
rect 10610 12010 10650 12050
rect 10690 12010 10730 12050
rect 10770 12010 10810 12050
rect 10850 12010 10890 12050
rect 10930 12010 10970 12050
rect 11010 12010 11050 12050
rect 11090 12010 11130 12050
rect 11170 12010 11210 12050
rect 11250 12010 11290 12050
rect 11330 12010 11370 12050
rect 11410 12010 11450 12050
rect 11490 12010 11530 12050
rect 11570 12010 11610 12050
rect 11650 12010 11690 12050
rect 11730 12010 11770 12050
rect 11810 12010 11850 12050
rect 11890 12010 11930 12050
rect 11970 12010 12010 12050
rect 12050 12010 12090 12050
rect 12130 12010 12170 12050
rect 12210 12010 12250 12050
rect 12290 12010 12330 12050
rect 12370 12010 12410 12050
rect 12450 12010 12490 12050
rect 12530 12010 12570 12050
rect 12610 12010 12650 12050
rect 12690 12010 12730 12050
rect 12770 12010 12810 12050
rect 12850 12010 12890 12050
rect 12930 12010 12970 12050
rect 13010 12010 13050 12050
rect 13090 12010 13130 12050
rect 13170 12010 13210 12050
rect 13250 12010 13290 12050
rect 13330 12010 13440 12050
rect 13480 12010 13520 12050
rect 13560 12010 13600 12050
rect 13640 12010 13680 12050
rect 13720 12010 13760 12050
rect 13800 12010 13840 12050
rect 13880 12010 13920 12050
rect 13960 12010 14000 12050
rect 14040 12010 14080 12050
rect 14120 12010 14160 12050
rect 14200 12010 14240 12050
rect 14280 12010 14320 12050
rect 14360 12010 14400 12050
rect 14440 12010 14480 12050
rect 14520 12010 14560 12050
rect 14600 12010 14640 12050
rect 14680 12010 14720 12050
rect 14760 12010 14800 12050
rect 14840 12010 14880 12050
rect 14920 12010 14960 12050
rect 15000 12010 15040 12050
rect 15080 12010 15120 12050
rect 15160 12010 15200 12050
rect 15240 12010 15280 12050
rect 15320 12010 15360 12050
rect 15400 12010 15440 12050
rect 15480 12010 15520 12050
rect 15560 12010 15600 12050
rect 15640 12010 15680 12050
rect 15720 12010 15760 12050
rect 15800 12010 15840 12050
rect 15880 12010 15920 12050
rect 15960 12010 16000 12050
rect 16040 12010 16080 12050
rect 16120 12010 16160 12050
rect 16200 12010 16240 12050
rect 16280 12010 16320 12050
rect 16360 12010 16400 12050
rect 16440 12010 16480 12050
rect 16520 12010 16560 12050
rect 16600 12010 16640 12050
rect 16680 12010 16720 12050
rect 16760 12010 16800 12050
rect 16840 12010 16880 12050
rect 16920 12010 16960 12050
rect 17000 12010 17040 12050
rect 17080 12010 17120 12050
rect 17160 12010 17200 12050
rect 17240 12010 17280 12050
rect 17320 12010 17360 12050
rect 17400 12010 17440 12050
rect 17480 12010 17520 12050
rect 17560 12010 17600 12050
rect 17640 12010 17680 12050
rect 17720 12010 17760 12050
rect 17800 12010 17840 12050
rect 17880 12010 17920 12050
rect 17960 12010 18000 12050
rect 18040 12010 18080 12050
rect 18120 12010 18160 12050
rect 18200 12010 18240 12050
rect 18280 12010 18320 12050
rect 18360 12010 18400 12050
rect 18440 12010 18480 12050
rect 18520 12010 18560 12050
rect 18600 12010 18640 12050
rect 18680 12010 18720 12050
rect 18760 12010 18800 12050
rect 18840 12010 18880 12050
rect 18920 12010 18960 12050
rect 19000 12010 19040 12050
rect 19080 12010 19120 12050
rect 19160 12010 19200 12050
rect 19240 12010 19280 12050
rect 19320 12010 19360 12050
rect 19400 12010 19440 12050
rect 19480 12010 19520 12050
rect 19560 12010 19600 12050
rect 19640 12010 19680 12050
rect 19720 12010 19760 12050
rect 19800 12010 19840 12050
rect 19890 12010 19930 12050
rect 19970 12010 20010 12050
rect 20050 12010 20090 12050
rect 20130 12010 20170 12050
rect 20210 12010 20250 12050
rect 20290 12010 20330 12050
rect 20370 12010 20410 12050
rect 20460 12010 20500 12050
rect 20540 12010 20580 12050
rect 20620 12010 20660 12050
rect 20700 12010 20740 12050
rect 20780 12010 20820 12050
rect 20860 12010 20900 12050
rect 20940 12010 20980 12050
rect 21020 12010 21060 12050
rect 7330 11960 7370 12000
rect 7410 11960 7450 12000
rect 7490 11960 7530 12000
rect 7570 11960 7610 12000
rect 7650 11960 7690 12000
rect 7730 11960 7770 12000
rect 7810 11960 7850 12000
rect 7890 11960 7930 12000
rect 7970 11960 8010 12000
rect 8050 11960 8090 12000
rect 8130 11960 8170 12000
rect 8210 11960 8250 12000
rect 8290 11960 8330 12000
rect 8370 11960 8410 12000
rect 8450 11960 8490 12000
rect 8530 11960 8570 12000
rect 8610 11960 8650 12000
rect 8690 11960 8730 12000
rect 8770 11960 8810 12000
rect 8850 11960 8890 12000
rect 8930 11960 8970 12000
rect 9010 11960 9050 12000
rect 9090 11960 9130 12000
rect 9170 11960 9210 12000
rect 9250 11960 9290 12000
rect 9330 11960 9370 12000
rect 9410 11960 9450 12000
rect 9490 11960 9530 12000
rect 9570 11960 9610 12000
rect 9650 11960 9690 12000
rect 9730 11960 9770 12000
rect 7720 11370 7760 11410
rect 7800 11370 7840 11410
rect 7880 11370 7920 11410
rect 7960 11370 8000 11410
rect 8040 11370 8080 11410
rect 8120 11370 8160 11410
rect 8200 11370 8240 11410
rect 8280 11370 8320 11410
rect 8360 11370 8400 11410
rect 8440 11370 8480 11410
rect 8520 11370 8560 11410
rect 7670 11290 7710 11330
rect 7670 11210 7710 11250
rect 7670 11130 7710 11170
rect 7330 11050 7370 11090
rect 7410 11050 7450 11090
rect 7490 11050 7530 11090
rect 7570 11050 7610 11090
rect 7650 11050 7690 11090
rect 7270 10350 7330 10410
rect 8550 11290 8590 11330
rect 8550 11210 8590 11250
rect 8550 11130 8590 11170
rect 8610 11050 8650 11090
rect 8690 11050 8730 11090
rect 8770 11050 8810 11090
rect 8850 11050 8890 11090
rect 8930 11050 8970 11090
rect 9010 11050 9050 11090
rect 9090 11050 9130 11090
rect 9170 11050 9210 11090
rect 9250 11050 9290 11090
rect 9330 11050 9370 11090
rect 9410 11050 9450 11090
rect 9490 11050 9530 11090
rect 9570 11050 9610 11090
rect 9650 11050 9690 11090
rect 9730 11050 9770 11090
rect 7610 10890 7670 10950
rect 8130 10900 8170 10940
rect 8350 10900 8390 10940
rect 7850 10790 7910 10850
rect 7610 10340 7650 10380
rect 7320 9680 7360 9720
rect 7400 9680 7440 9720
rect 7480 9680 7520 9720
rect 7560 9680 7600 9720
rect 7640 9680 7680 9720
rect 7720 9680 7760 9720
rect 8810 10480 8850 10520
rect 9810 11000 9850 11040
rect 9890 11000 9930 11040
rect 9970 11000 10010 11040
rect 10050 11000 10090 11040
rect 10130 11000 10170 11040
rect 10210 11000 10250 11040
rect 10290 11000 10330 11040
rect 10370 11000 10410 11040
rect 10450 11000 10490 11040
rect 10530 11000 10570 11040
rect 10610 11000 10650 11040
rect 10690 11000 10730 11040
rect 10770 11000 10810 11040
rect 10850 11000 10890 11040
rect 10930 11000 10970 11040
rect 11010 11000 11050 11040
rect 11090 11000 11130 11040
rect 11170 11000 11210 11040
rect 11250 11000 11290 11040
rect 11330 11000 11370 11040
rect 11410 11000 11450 11040
rect 11490 11000 11530 11040
rect 11570 11000 11610 11040
rect 11650 11000 11690 11040
rect 11730 11000 11770 11040
rect 11810 11000 11850 11040
rect 11890 11000 11930 11040
rect 11970 11000 12010 11040
rect 12050 11000 12090 11040
rect 12130 11000 12170 11040
rect 12210 11000 12250 11040
rect 12290 11000 12330 11040
rect 12370 11000 12410 11040
rect 12450 11000 12490 11040
rect 12530 11000 12570 11040
rect 12610 11000 12650 11040
rect 12690 11000 12730 11040
rect 12770 11000 12810 11040
rect 12850 11000 12890 11040
rect 12930 11000 12970 11040
rect 13010 11000 13050 11040
rect 13090 11000 13130 11040
rect 13170 11000 13210 11040
rect 13250 11000 13290 11040
rect 13330 11000 13410 11040
rect 13450 11000 13490 11040
rect 13530 11000 13570 11040
rect 13610 11000 13650 11040
rect 13690 11000 13730 11040
rect 13770 11000 13810 11040
rect 13850 11000 13890 11040
rect 13930 11000 13970 11040
rect 14010 11000 14050 11040
rect 14090 11000 14130 11040
rect 14170 11000 14210 11040
rect 14250 11000 14290 11040
rect 14330 11000 14370 11040
rect 14410 11000 14450 11040
rect 14490 11000 14530 11040
rect 14570 11000 14610 11040
rect 14650 11000 14690 11040
rect 14730 11000 14770 11040
rect 14810 11000 14850 11040
rect 14890 11000 14930 11040
rect 14970 11000 15010 11040
rect 15050 11000 15090 11040
rect 15130 11000 15170 11040
rect 15210 11000 15250 11040
rect 15290 11000 15330 11040
rect 15370 11000 15410 11040
rect 15450 11000 15490 11040
rect 15530 11000 15570 11040
rect 15610 11000 15650 11040
rect 15690 11000 15730 11040
rect 15770 11000 15810 11040
rect 15850 11000 15890 11040
rect 15930 11000 15970 11040
rect 16010 11000 16050 11040
rect 16090 11000 16130 11040
rect 16170 11000 16210 11040
rect 16250 11000 16290 11040
rect 16330 11000 16370 11040
rect 16410 11000 16450 11040
rect 16490 11000 16530 11040
rect 16570 11000 16610 11040
rect 16650 11000 16690 11040
rect 16730 11000 16770 11040
rect 16810 11000 16850 11040
rect 16890 11000 16930 11040
rect 16970 11000 17010 11040
rect 17050 11000 17090 11040
rect 17130 11000 17170 11040
rect 17210 11000 17250 11040
rect 17290 11000 17330 11040
rect 17370 11000 17410 11040
rect 17450 11000 17490 11040
rect 17530 11000 17570 11040
rect 17610 11000 17650 11040
rect 17690 11000 17730 11040
rect 17770 11000 17810 11040
rect 17850 11000 17890 11040
rect 17930 11000 17970 11040
rect 18010 11000 18050 11040
rect 18090 11000 18130 11040
rect 18170 11000 18210 11040
rect 18250 11000 18290 11040
rect 18330 11000 18370 11040
rect 18410 11000 18450 11040
rect 18490 11000 18530 11040
rect 18570 11000 18610 11040
rect 18650 11000 18690 11040
rect 18730 11000 18770 11040
rect 18810 11000 18850 11040
rect 18890 11000 18930 11040
rect 18970 11000 19010 11040
rect 19050 11000 19090 11040
rect 19130 11000 19170 11040
rect 19210 11000 19250 11040
rect 19290 11000 19330 11040
rect 19370 11000 19410 11040
rect 19450 11000 19490 11040
rect 19540 11000 19580 11040
rect 19620 11000 19660 11040
rect 19700 11000 19740 11040
rect 19780 11000 19820 11040
rect 19860 11000 19900 11040
rect 19940 11000 19980 11040
rect 20020 11000 20060 11040
rect 20110 11000 20150 11040
rect 20190 11000 20230 11040
rect 20270 11000 20310 11040
rect 20350 11000 20390 11040
rect 20430 11000 20470 11040
rect 20510 11000 20550 11040
rect 20590 11000 20630 11040
rect 20670 11000 20710 11040
rect 20750 11000 20790 11040
rect 20830 11000 20870 11040
rect 20910 11000 20950 11040
rect 20990 11000 21030 11040
rect 21070 11000 21110 11040
rect 9650 10780 9720 10840
rect 9860 10640 9900 10680
rect 8660 10370 8700 10410
rect 8960 10360 9000 10400
rect 9040 10360 9080 10400
rect 9160 10360 9200 10400
rect 9300 10360 9340 10400
rect 9420 10360 9460 10400
rect 9550 10360 9590 10400
rect 9670 10360 9710 10400
rect 9790 10350 9860 10410
rect 10680 10450 10720 10490
rect 11290 10470 11360 10530
rect 11670 10450 11710 10490
rect 12290 10440 12360 10500
rect 12670 10450 12710 10490
rect 10160 10340 10200 10380
rect 10420 10350 10460 10390
rect 10920 10340 10960 10380
rect 11000 10340 11040 10380
rect 11300 10340 11340 10380
rect 11410 10350 11450 10390
rect 11910 10340 11950 10380
rect 11990 10340 12030 10380
rect 12290 10340 12330 10380
rect 12410 10350 12450 10390
rect 12910 10340 12950 10380
rect 12990 10340 13030 10380
rect 13270 10350 13310 10390
rect 13350 10350 13390 10390
rect 13450 10350 13490 10390
rect 13580 10350 13620 10390
rect 13790 10350 13830 10390
rect 13920 10350 13960 10390
rect 14350 10350 14390 10390
rect 14480 10350 14520 10390
rect 15350 10350 15390 10390
rect 15540 10350 15580 10390
rect 17340 10350 17390 10400
rect 17490 10350 17530 10390
rect 21050 10350 21100 10400
rect 8520 9680 8560 9720
rect 8600 9680 8640 9720
rect 8680 9680 8720 9720
rect 8760 9680 8800 9720
rect 8840 9680 8880 9720
rect 8920 9680 8960 9720
rect 9000 9680 9040 9720
rect 9080 9680 9120 9720
rect 9160 9680 9200 9720
rect 9240 9680 9280 9720
rect 9320 9680 9360 9720
rect 9400 9680 9440 9720
rect 9480 9680 9520 9720
rect 9560 9680 9600 9720
rect 9640 9680 9680 9720
rect 9720 9680 9760 9720
rect 9800 9680 9840 9720
rect 9890 9680 9930 9720
rect 9970 9680 10010 9720
rect 10050 9680 10090 9720
rect 10130 9680 10170 9720
rect 10210 9680 10250 9720
rect 10290 9680 10330 9720
rect 10370 9680 10410 9720
rect 10450 9680 10490 9720
rect 10530 9680 10570 9720
rect 10610 9680 10650 9720
rect 10690 9680 10730 9720
rect 10770 9680 10810 9720
rect 10850 9680 10890 9720
rect 10930 9680 10970 9720
rect 11010 9680 11050 9720
rect 11090 9680 11130 9720
rect 11170 9680 11210 9720
rect 11250 9680 11290 9720
rect 11330 9680 11370 9720
rect 11410 9680 11450 9720
rect 11490 9680 11530 9720
rect 11570 9680 11610 9720
rect 11650 9680 11690 9720
rect 11730 9680 11770 9720
rect 11810 9680 11850 9720
rect 11890 9680 11930 9720
rect 11970 9680 12010 9720
rect 12050 9680 12090 9720
rect 12130 9680 12170 9720
rect 12210 9680 12250 9720
rect 12290 9680 12330 9720
rect 12370 9680 12410 9720
rect 12450 9680 12490 9720
rect 12530 9680 12570 9720
rect 12610 9680 12650 9720
rect 12690 9680 12730 9720
rect 12770 9680 12810 9720
rect 12850 9680 12890 9720
rect 12930 9680 12970 9720
rect 13010 9680 13050 9720
rect 13090 9680 13130 9720
rect 13170 9680 13210 9720
rect 13250 9680 13290 9720
rect 13330 9680 13370 9720
rect 13410 9680 13450 9720
rect 13490 9680 13530 9720
rect 13570 9680 13610 9720
rect 13650 9680 13690 9720
rect 13730 9680 13770 9720
rect 13810 9680 13850 9720
rect 13890 9680 13930 9720
rect 13970 9680 14010 9720
rect 14050 9680 14090 9720
rect 14130 9680 14170 9720
rect 14210 9680 14250 9720
rect 14290 9680 14330 9720
rect 14370 9680 14410 9720
rect 14450 9680 14490 9720
rect 14530 9680 14570 9720
rect 14610 9680 14650 9720
rect 14690 9680 14730 9720
rect 14770 9680 14810 9720
rect 14850 9680 14890 9720
rect 14930 9680 14970 9720
rect 15010 9680 15050 9720
rect 15090 9680 15130 9720
rect 15170 9680 15210 9720
rect 15250 9680 15290 9720
rect 15330 9680 15370 9720
rect 15410 9680 15450 9720
rect 15490 9680 15530 9720
rect 15570 9680 15610 9720
rect 15650 9680 15690 9720
rect 15730 9680 15770 9720
rect 15810 9680 15850 9720
rect 15890 9680 15930 9720
rect 15970 9680 16010 9720
rect 16050 9680 16090 9720
rect 16130 9680 16170 9720
rect 16210 9680 16250 9720
rect 16290 9680 16330 9720
rect 16370 9680 16410 9720
rect 16450 9680 16490 9720
rect 16530 9680 16570 9720
rect 16610 9680 16650 9720
rect 16690 9680 16730 9720
rect 16770 9680 16810 9720
rect 16850 9680 16890 9720
rect 16930 9680 16970 9720
rect 17010 9680 17050 9720
rect 17090 9680 17130 9720
rect 17170 9680 17210 9720
rect 17250 9680 17290 9720
rect 17330 9680 17370 9720
rect 17410 9680 17450 9720
rect 17490 9680 17530 9720
rect 17570 9680 17610 9720
rect 17650 9680 17690 9720
rect 17730 9680 17770 9720
rect 17810 9680 17850 9720
rect 17890 9680 17930 9720
rect 17970 9680 18010 9720
rect 18050 9680 18090 9720
rect 18130 9680 18170 9720
rect 18210 9680 18250 9720
rect 18290 9680 18330 9720
rect 18370 9680 18410 9720
rect 18450 9680 18490 9720
rect 18530 9680 18570 9720
rect 18610 9680 18650 9720
rect 18690 9680 18730 9720
rect 18770 9680 18810 9720
rect 18850 9680 18890 9720
rect 18930 9680 18970 9720
rect 19010 9680 19050 9720
rect 19090 9680 19130 9720
rect 19170 9680 19210 9720
rect 19250 9680 19290 9720
rect 19330 9680 19370 9720
rect 19410 9680 19450 9720
rect 19490 9680 19530 9720
rect 19570 9680 19610 9720
rect 19650 9680 19690 9720
rect 19730 9680 19770 9720
rect 19810 9680 19850 9720
rect 19890 9680 19930 9720
rect 19970 9680 20010 9720
rect 20050 9680 20090 9720
rect 20130 9680 20170 9720
rect 20210 9680 20250 9720
rect 20290 9680 20330 9720
rect 20370 9680 20410 9720
rect 20450 9680 20490 9720
rect 20530 9680 20570 9720
rect 20610 9680 20650 9720
rect 20690 9680 20730 9720
rect 20770 9680 20810 9720
rect 20850 9680 20890 9720
rect 20930 9680 20970 9720
rect 21010 9680 21050 9720
rect 7740 9590 7780 9630
rect 7820 9590 7860 9630
rect 7900 9590 7940 9630
rect 7980 9590 8020 9630
rect 8060 9590 8100 9630
rect 8140 9590 8180 9630
rect 8220 9590 8260 9630
rect 8300 9590 8340 9630
rect 8380 9590 8420 9630
rect 8460 9590 8500 9630
rect 21570 8850 21640 8920
rect 21970 8850 22040 8920
rect 22400 8850 22470 8920
rect 13220 8580 13270 8630
rect 22570 8570 22640 8640
rect 23270 8570 23340 8640
rect 13430 8420 13560 8490
rect 17050 8310 17100 8360
rect 9900 6930 9960 6980
rect 10120 6930 10180 6980
rect 10340 6930 10400 6980
rect 10560 6930 10620 6980
rect 10780 6930 10840 6980
rect 11000 6930 11060 6980
rect 11220 6930 11280 6980
rect 11440 6930 11500 6980
rect 11660 6930 11720 6980
rect 11880 6930 11940 6980
rect 12100 6930 12160 6980
rect 12320 6930 12380 6980
rect 12540 6930 12600 6980
rect 12760 6930 12820 6980
rect 12980 6930 13040 6980
rect 13200 6930 13260 6980
rect 13670 6930 13730 6980
rect 13890 6930 13950 6980
rect 14110 6930 14170 6980
rect 14330 6930 14390 6980
rect 14550 6930 14610 6980
rect 14770 6930 14830 6980
rect 14990 6930 15050 6980
rect 15210 6930 15270 6980
rect 15430 6930 15490 6980
rect 15650 6930 15710 6980
rect 15870 6930 15930 6980
rect 16090 6930 16150 6980
rect 16310 6930 16370 6980
rect 16530 6930 16590 6980
rect 16750 6930 16810 6980
rect 16970 6930 17030 6980
rect 13630 5940 13690 5990
rect 13850 5940 13910 5990
rect 14070 5940 14130 5990
rect 14290 5940 14350 5990
rect 14510 5940 14570 5990
rect 14730 5940 14790 5990
rect 14950 5940 15010 5990
rect 15170 5940 15230 5990
rect 15390 5940 15450 5990
rect 15610 5940 15670 5990
rect 15830 5940 15890 5990
rect 16050 5940 16110 5990
rect 16270 5940 16330 5990
rect 16490 5940 16550 5990
rect 16710 5940 16770 5990
rect 16930 5940 16990 5990
rect 9930 5830 9970 5870
rect 10010 5830 10050 5870
rect 10090 5830 10130 5870
rect 10170 5830 10210 5870
rect 10250 5830 10290 5870
rect 10330 5830 10370 5870
rect 10410 5830 10450 5870
rect 10490 5830 10530 5870
rect 10610 5830 10650 5870
rect 10690 5830 10730 5870
rect 10770 5830 10810 5870
rect 10850 5830 10890 5870
rect 10930 5830 10970 5870
rect 11010 5830 11050 5870
rect 11090 5830 11130 5870
rect 11170 5830 11210 5870
rect 11250 5830 11290 5870
rect 11370 5830 11410 5870
rect 11450 5830 11490 5870
rect 11530 5830 11570 5870
rect 11610 5830 11650 5870
rect 11690 5830 11730 5870
rect 11770 5830 11810 5870
rect 11850 5830 11890 5870
rect 11930 5830 11970 5870
rect 12010 5830 12050 5870
rect 12130 5830 12170 5870
rect 12210 5830 12250 5870
rect 12290 5830 12330 5870
rect 12370 5830 12410 5870
rect 12450 5830 12490 5870
rect 12530 5830 12570 5870
rect 12610 5830 12650 5870
rect 12690 5830 12730 5870
rect 12770 5830 12810 5870
rect 12850 5830 12890 5870
rect 12930 5830 12970 5870
rect 13010 5830 13050 5870
rect 13090 5830 13130 5870
rect 13380 5820 13510 5880
rect 9850 4070 9930 4140
rect 13380 4440 13510 4500
rect 16950 4420 17000 4470
rect 13380 4280 13510 4340
rect 13180 4090 13250 4150
rect 13180 3900 13250 3960
rect 21970 4240 22040 4310
rect 22400 4240 22470 4310
rect 13320 3020 13450 3080
rect 16950 3190 17000 3240
rect 13630 2950 13690 3000
rect 13850 2950 13910 3000
rect 14070 2950 14130 3000
rect 14290 2950 14350 3000
rect 14510 2950 14570 3000
rect 14730 2950 14790 3000
rect 14950 2950 15010 3000
rect 15170 2950 15230 3000
rect 15390 2950 15450 3000
rect 15610 2950 15670 3000
rect 15830 2950 15890 3000
rect 16050 2950 16110 3000
rect 16270 2950 16330 3000
rect 16490 2950 16550 3000
rect 16710 2950 16770 3000
rect 24220 2660 24280 2720
rect 24220 2560 24280 2620
rect 25720 2720 25770 2760
rect 25720 2600 25770 2640
rect 24220 2460 24280 2520
rect 24220 2360 24280 2420
rect 25720 2480 25770 2520
rect 25720 2360 25770 2400
rect 24220 2260 24280 2320
rect 24220 2160 24280 2220
rect 24220 2060 24280 2120
rect 25720 2240 25770 2280
rect 25720 2120 25770 2160
rect 9890 1870 9950 1920
rect 10110 1870 10170 1920
rect 10330 1870 10390 1920
rect 10550 1870 10610 1920
rect 10770 1870 10830 1920
rect 10990 1870 11050 1920
rect 11210 1870 11270 1920
rect 11430 1870 11490 1920
rect 11650 1870 11710 1920
rect 11870 1870 11930 1920
rect 12090 1870 12150 1920
rect 12310 1870 12370 1920
rect 12530 1870 12590 1920
rect 12750 1870 12810 1920
rect 12970 1870 13030 1920
rect 13630 1870 13690 1920
rect 13850 1870 13910 1920
rect 14070 1870 14130 1920
rect 14290 1870 14350 1920
rect 14510 1870 14570 1920
rect 14730 1870 14790 1920
rect 14950 1870 15010 1920
rect 15170 1870 15230 1920
rect 15390 1870 15450 1920
rect 15610 1870 15670 1920
rect 15830 1870 15890 1920
rect 16050 1870 16110 1920
rect 16270 1870 16330 1920
rect 16490 1870 16550 1920
rect 16710 1870 16770 1920
rect 25480 1910 25540 1970
rect 13210 1630 13260 1680
rect 13360 530 13490 600
rect 17060 1370 17110 1420
rect 21570 350 21640 420
<< metal1 >>
rect 2070 44100 3000 44160
rect 2070 43410 2120 44100
rect 2950 43410 3000 44100
rect 2070 42170 3000 43410
rect 21680 44100 23880 44160
rect 21680 43410 21730 44100
rect 22580 43410 22980 44100
rect 23830 43410 23880 44100
rect 21680 43360 23880 43410
rect 21790 43350 23880 43360
rect 21790 43280 21830 43350
rect 21890 43280 21930 43350
rect 21990 43280 22030 43350
rect 22090 43280 22130 43350
rect 22190 43280 22230 43350
rect 22290 43280 22330 43350
rect 22390 43280 22430 43350
rect 22490 43280 22530 43350
rect 22590 43280 22630 43350
rect 22690 43280 22730 43350
rect 22790 43280 22830 43350
rect 22890 43280 22930 43350
rect 22990 43280 23030 43350
rect 23090 43280 23130 43350
rect 23190 43280 23230 43350
rect 23290 43280 23330 43350
rect 23390 43280 23430 43350
rect 23490 43280 23530 43350
rect 23590 43280 23880 43350
rect 21790 43270 23880 43280
rect 15670 43180 15790 43200
rect 3380 43000 4330 43060
rect 15670 43050 15690 43180
rect 15770 43050 15790 43180
rect 22320 43150 22420 43170
rect 22320 43090 22340 43150
rect 22400 43090 22420 43150
rect 22320 43070 22420 43090
rect 15670 43030 15790 43050
rect 3380 42310 3430 43000
rect 4280 42310 4330 43000
rect 3380 42260 4330 42310
rect 2439 42160 3159 42170
rect 2439 42110 2469 42160
rect 2519 42110 2559 42160
rect 2609 42110 2649 42160
rect 2699 42110 2739 42160
rect 2789 42110 2829 42160
rect 2879 42110 2919 42160
rect 2969 42110 3159 42160
rect 2439 42100 3159 42110
rect 2769 42050 2849 42060
rect 2769 42010 2789 42050
rect 2829 42010 2849 42050
rect 2769 42000 2849 42010
rect 3099 41800 3159 42100
rect 3380 41950 4329 42260
rect 5619 41980 9979 42040
rect 3380 41900 3429 41950
rect 3479 41900 3519 41950
rect 3569 41900 3609 41950
rect 3659 41900 3699 41950
rect 3749 41900 3789 41950
rect 3839 41900 3879 41950
rect 3929 41900 3969 41950
rect 4019 41900 4059 41950
rect 4109 41900 4149 41950
rect 4199 41900 4239 41950
rect 4289 41900 4329 41950
rect 3380 41890 4329 41900
rect 4539 41950 5479 41960
rect 4539 41890 4579 41950
rect 4639 41890 5479 41950
rect 4539 41880 5479 41890
rect 3099 41750 3340 41800
rect 3049 41690 3209 41700
rect 3049 41630 3079 41690
rect 3179 41630 3209 41690
rect 2659 41620 2739 41630
rect 3049 41620 3209 41630
rect 2659 41580 2679 41620
rect 2719 41580 2739 41620
rect 2659 41570 2739 41580
rect 2879 41580 2959 41590
rect 3089 41580 3129 41620
rect 2879 41540 2899 41580
rect 2939 41540 3129 41580
rect 2879 41530 2959 41540
rect 2779 41510 2839 41530
rect 2779 41470 2789 41510
rect 2829 41500 2839 41510
rect 3159 41520 3259 41530
rect 3159 41500 3179 41520
rect 2829 41470 3179 41500
rect 2779 41450 2839 41470
rect 3159 41460 3179 41470
rect 3239 41460 3259 41520
rect 3159 41450 3259 41460
rect 3290 40990 3340 41750
rect 3459 40990 3519 41010
rect 2979 40940 3039 40960
rect 3290 40950 3469 40990
rect 3509 40950 3519 40990
rect 2979 40900 2989 40940
rect 3029 40900 3039 40940
rect 3459 40930 3519 40950
rect 5349 40980 5409 41000
rect 5349 40940 5359 40980
rect 5399 40940 5409 40980
rect 5349 40920 5409 40940
rect 5489 40920 5589 40930
rect 2979 40880 3039 40900
rect 5489 40860 5509 40920
rect 5569 40910 5589 40920
rect 5619 40910 5689 41980
rect 5939 41970 9979 41980
rect 5939 41910 6009 41970
rect 6069 41910 6119 41970
rect 6179 41910 6229 41970
rect 6289 41910 6339 41970
rect 6399 41910 6449 41970
rect 6509 41910 6559 41970
rect 6619 41910 6669 41970
rect 6729 41910 6779 41970
rect 6839 41910 6889 41970
rect 6949 41910 6999 41970
rect 7059 41910 7109 41970
rect 7169 41910 7219 41970
rect 7279 41910 7329 41970
rect 7389 41910 7439 41970
rect 7499 41910 7549 41970
rect 7609 41910 7659 41970
rect 7719 41910 7769 41970
rect 7829 41910 7879 41970
rect 7939 41910 7989 41970
rect 8049 41910 8099 41970
rect 8159 41910 8209 41970
rect 8269 41910 8319 41970
rect 8379 41910 8429 41970
rect 8489 41910 8539 41970
rect 8599 41910 8649 41970
rect 8709 41910 8759 41970
rect 8819 41910 8869 41970
rect 8929 41910 8979 41970
rect 9039 41910 9089 41970
rect 9149 41910 9199 41970
rect 9259 41910 9309 41970
rect 9369 41910 9419 41970
rect 9479 41910 9529 41970
rect 9589 41910 9639 41970
rect 9699 41910 9749 41970
rect 9809 41910 9859 41970
rect 9919 41910 9979 41970
rect 5939 41900 9979 41910
rect 15690 42000 15770 43030
rect 22220 42960 23260 43000
rect 22050 42130 22150 42140
rect 22050 42070 22070 42130
rect 22130 42070 22150 42130
rect 22050 42060 22150 42070
rect 15690 41980 21780 42000
rect 15690 41920 21630 41980
rect 21700 41920 21780 41980
rect 21820 41970 21910 41980
rect 22220 41970 22260 42960
rect 23220 42320 23260 42960
rect 23450 42320 23530 42330
rect 23220 42280 23470 42320
rect 23510 42280 23530 42320
rect 23450 42270 23530 42280
rect 23800 42220 23880 43270
rect 23480 42210 23880 42220
rect 23480 42170 23500 42210
rect 23540 42170 23880 42210
rect 23480 42160 23880 42170
rect 23090 42140 23170 42150
rect 22570 42100 22650 42110
rect 22570 42060 22590 42100
rect 22630 42060 22650 42100
rect 23090 42100 23110 42140
rect 23150 42100 23170 42140
rect 23090 42090 23170 42100
rect 22570 42050 22650 42060
rect 22580 41990 22630 42050
rect 22980 42030 23060 42040
rect 23110 42030 23150 42090
rect 22980 41990 23000 42030
rect 23040 41990 23150 42030
rect 22580 41970 22650 41990
rect 22980 41980 23060 41990
rect 21820 41930 21850 41970
rect 21890 41930 22590 41970
rect 22630 41930 22650 41970
rect 21820 41920 21910 41930
rect 15690 41900 21780 41920
rect 22580 41910 22650 41930
rect 23110 41970 23190 41990
rect 23110 41930 23120 41970
rect 23160 41930 23190 41970
rect 22980 41910 23060 41920
rect 23110 41910 23190 41930
rect 22580 41810 22630 41910
rect 22980 41870 23000 41910
rect 23040 41870 23150 41910
rect 22980 41860 23060 41870
rect 23110 41810 23150 41870
rect 23620 41870 23740 41890
rect 23620 41810 23640 41870
rect 23720 41810 23740 41870
rect 22570 41800 22650 41810
rect 22570 41760 22590 41800
rect 22630 41760 22650 41800
rect 22570 41750 22650 41760
rect 23090 41800 23170 41810
rect 23090 41760 23110 41800
rect 23150 41760 23170 41800
rect 23620 41790 23740 41810
rect 23090 41750 23170 41760
rect 23480 41760 23560 41770
rect 23480 41720 23500 41760
rect 23540 41720 23560 41760
rect 23480 41710 23560 41720
rect 23800 41690 23880 42160
rect 23800 41630 23810 41690
rect 23870 41630 23880 41690
rect 23800 41610 23880 41630
rect 22430 41330 22530 41350
rect 5959 41280 6019 41300
rect 5569 40870 5689 40910
rect 5719 41240 5969 41280
rect 6009 41240 6019 41280
rect 5569 40860 5589 40870
rect 5489 40850 5589 40860
rect 5719 40790 5759 41240
rect 5959 41220 6019 41240
rect 6059 41280 6249 41300
rect 6059 41240 6069 41280
rect 6109 41240 6199 41280
rect 6239 41240 6249 41280
rect 6059 41220 6249 41240
rect 6399 41280 6589 41300
rect 6399 41240 6409 41280
rect 6449 41240 6539 41280
rect 6579 41240 6589 41280
rect 6399 41220 6589 41240
rect 6959 41280 7149 41300
rect 6959 41240 6969 41280
rect 7009 41240 7099 41280
rect 7139 41240 7149 41280
rect 6959 41220 7149 41240
rect 7959 41280 8209 41300
rect 7959 41240 7969 41280
rect 8009 41240 8159 41280
rect 8199 41240 8209 41280
rect 7959 41220 8209 41240
rect 9899 41280 10029 41290
rect 9899 41230 9959 41280
rect 10009 41230 10119 41280
rect 22430 41270 22450 41330
rect 22510 41270 22530 41330
rect 22430 41250 22530 41270
rect 9899 41220 10029 41230
rect 5949 40910 9979 40920
rect 5949 40850 6009 40910
rect 6070 40850 9979 40910
rect 5949 40840 9979 40850
rect 2869 40780 5759 40790
rect 2869 40770 3099 40780
rect 2869 40730 2879 40770
rect 2919 40740 3099 40770
rect 3139 40740 4419 40780
rect 4459 40740 5459 40780
rect 5499 40740 5759 40780
rect 2919 40730 5759 40740
rect 2869 40710 2929 40730
rect 2759 40660 3049 40680
rect 2759 40620 2769 40660
rect 2809 40620 2999 40660
rect 3039 40620 3049 40660
rect 2759 40600 3049 40620
rect 3260 40670 4200 40680
rect 3260 40610 3320 40670
rect 3380 40610 3430 40670
rect 3490 40610 3540 40670
rect 3600 40610 3650 40670
rect 3710 40610 3760 40670
rect 3820 40610 3870 40670
rect 3930 40610 3980 40670
rect 4040 40610 4090 40670
rect 4150 40610 4200 40670
rect 3260 40600 4200 40610
rect 4539 40660 5429 40680
rect 4539 40620 4659 40660
rect 5399 40620 5429 40660
rect 4539 40600 5429 40620
rect 2869 40530 2929 40550
rect 2869 40490 2879 40530
rect 2919 40490 2929 40530
rect 2749 39690 2809 39710
rect 2869 39690 2929 40490
rect 2749 39650 2759 39690
rect 2799 39650 2929 39690
rect 3329 39700 3389 39720
rect 3329 39660 3339 39700
rect 3379 39660 3389 39700
rect 2749 39630 2809 39650
rect 2070 39570 2620 39580
rect 3329 39570 3389 39660
rect 5349 39700 5409 39720
rect 5349 39660 5359 39700
rect 5399 39660 5409 39700
rect 5349 39570 5409 39660
rect 6009 39570 6069 40840
rect 10069 40750 10119 41230
rect 21590 41160 23630 41180
rect 21590 41090 21620 41160
rect 21680 41090 21720 41160
rect 21780 41090 21830 41160
rect 21890 41090 21930 41160
rect 21990 41090 22030 41160
rect 22090 41090 22130 41160
rect 22190 41090 22230 41160
rect 22290 41090 22330 41160
rect 22390 41090 22430 41160
rect 22490 41090 22530 41160
rect 22590 41090 22630 41160
rect 22690 41090 22730 41160
rect 22790 41090 22830 41160
rect 22890 41090 22930 41160
rect 22990 41090 23030 41160
rect 23090 41090 23130 41160
rect 23190 41090 23230 41160
rect 23290 41090 23330 41160
rect 23390 41090 23430 41160
rect 23490 41090 23530 41160
rect 23590 41090 23630 41160
rect 21590 41080 23630 41090
rect 6179 40700 10119 40750
rect 21560 41020 23950 41080
rect 6179 39960 6219 40700
rect 6349 40650 9969 40660
rect 6349 40590 6409 40650
rect 6469 40590 6519 40650
rect 6579 40590 6629 40650
rect 6689 40590 6739 40650
rect 6799 40590 6849 40650
rect 6909 40590 6959 40650
rect 7019 40590 7069 40650
rect 7129 40590 7179 40650
rect 7239 40590 7289 40650
rect 7349 40590 7399 40650
rect 7459 40590 7509 40650
rect 7569 40590 7619 40650
rect 7679 40590 7729 40650
rect 7789 40590 7839 40650
rect 7899 40590 7949 40650
rect 8009 40590 8059 40650
rect 8119 40590 8169 40650
rect 8229 40590 8279 40650
rect 8339 40590 8389 40650
rect 8449 40590 8499 40650
rect 8559 40590 8609 40650
rect 8669 40590 8719 40650
rect 8779 40590 8829 40650
rect 8889 40590 8939 40650
rect 8999 40590 9049 40650
rect 9109 40590 9159 40650
rect 9219 40590 9269 40650
rect 9329 40590 9379 40650
rect 9439 40590 9489 40650
rect 9549 40590 9599 40650
rect 9659 40590 9709 40650
rect 9769 40590 9819 40650
rect 9879 40590 9969 40650
rect 6349 40580 9969 40590
rect 21560 40340 21610 41020
rect 22250 40340 22440 41020
rect 23080 40340 23260 41020
rect 23900 40340 23950 41020
rect 21560 40290 23950 40340
rect 10030 40000 10930 40020
rect 6349 39960 6419 39980
rect 10030 39970 10060 40000
rect 6179 39920 6369 39960
rect 6409 39920 6419 39960
rect 6349 39900 6419 39920
rect 9869 39960 10060 39970
rect 9869 39910 9929 39960
rect 9979 39910 10060 39960
rect 9869 39900 10060 39910
rect 10030 39880 10060 39900
rect 10900 39880 10930 40000
rect 10030 39860 10930 39880
rect 2070 39560 9979 39570
rect 2070 39500 2649 39560
rect 2709 39500 2749 39560
rect 2809 39500 2849 39560
rect 2909 39500 2949 39560
rect 3009 39500 3049 39560
rect 3109 39500 3149 39560
rect 3209 39500 3249 39560
rect 3309 39500 3349 39560
rect 3409 39500 3449 39560
rect 3509 39500 3549 39560
rect 3609 39500 3649 39560
rect 3709 39500 3749 39560
rect 3809 39500 3849 39560
rect 3909 39500 3949 39560
rect 4009 39500 4049 39560
rect 4109 39500 4149 39560
rect 4209 39500 4249 39560
rect 4309 39500 4349 39560
rect 4409 39500 4449 39560
rect 4509 39500 4549 39560
rect 4609 39500 4649 39560
rect 4709 39500 4749 39560
rect 4809 39500 4849 39560
rect 4909 39500 4949 39560
rect 5009 39500 5049 39560
rect 5109 39500 5149 39560
rect 5209 39500 5249 39560
rect 5309 39500 6349 39560
rect 6409 39500 6449 39560
rect 6509 39500 6549 39560
rect 6609 39500 6649 39560
rect 6709 39500 6749 39560
rect 6809 39500 6849 39560
rect 6909 39500 6949 39560
rect 7009 39500 7049 39560
rect 7109 39500 7149 39560
rect 7209 39500 7249 39560
rect 7309 39500 7349 39560
rect 7409 39500 7479 39560
rect 7539 39500 7579 39560
rect 7639 39500 7679 39560
rect 7739 39500 7779 39560
rect 7839 39500 7879 39560
rect 7939 39500 7979 39560
rect 8039 39500 8079 39560
rect 8139 39500 8179 39560
rect 8239 39500 8279 39560
rect 8339 39500 8379 39560
rect 8439 39500 8479 39560
rect 8539 39500 8629 39560
rect 8689 39500 8729 39560
rect 8789 39500 8829 39560
rect 8889 39500 8929 39560
rect 8989 39500 9029 39560
rect 9089 39500 9129 39560
rect 9189 39500 9229 39560
rect 9289 39500 9329 39560
rect 9389 39500 9429 39560
rect 9489 39500 9529 39560
rect 9589 39500 9629 39560
rect 9689 39500 9739 39560
rect 9799 39500 9839 39560
rect 9899 39500 9979 39560
rect 2070 39490 9979 39500
rect 2070 39430 9980 39490
rect 2070 38620 2130 39430
rect 3170 38620 3380 39430
rect 4420 38620 4630 39430
rect 5670 38620 5880 39430
rect 6920 38620 7130 39430
rect 8170 38620 8380 39430
rect 9850 38620 9980 39430
rect 2070 38560 9980 38620
rect 25320 38510 25410 38520
rect 25830 38510 25920 38520
rect 25320 38500 25920 38510
rect 25320 38430 25330 38500
rect 25400 38430 25840 38500
rect 25910 38430 25920 38500
rect 25320 38420 25920 38430
rect 25320 38410 25410 38420
rect 25830 38410 25920 38420
rect 2070 38050 10930 38110
rect 2070 37240 2120 38050
rect 3860 37240 4070 38050
rect 5110 37240 5320 38050
rect 6360 37240 6570 38050
rect 7610 37240 7820 38050
rect 8860 37240 9070 38050
rect 9820 37240 10080 38050
rect 10880 37240 10930 38050
rect 2070 37180 10930 37240
rect 2070 37120 3810 37180
rect 3870 37120 3910 37180
rect 3970 37120 4010 37180
rect 4070 37120 4110 37180
rect 4170 37120 4210 37180
rect 4270 37120 4310 37180
rect 4370 37120 4410 37180
rect 4470 37120 4510 37180
rect 4570 37120 4610 37180
rect 4670 37120 4710 37180
rect 4770 37120 4810 37180
rect 4870 37120 4910 37180
rect 4970 37120 5010 37180
rect 5070 37120 5110 37180
rect 5170 37120 5210 37180
rect 5270 37120 5310 37180
rect 5370 37120 5410 37180
rect 5470 37120 5510 37180
rect 5570 37120 5610 37180
rect 5670 37120 5710 37180
rect 5770 37120 5810 37180
rect 5870 37120 5910 37180
rect 5970 37120 6010 37180
rect 6070 37120 6110 37180
rect 6170 37120 10930 37180
rect 2070 37110 10930 37120
rect 2070 37100 3770 37110
rect 6340 36720 10930 37110
rect 6340 36660 6380 36720
rect 6440 36660 6480 36720
rect 6540 36660 6580 36720
rect 6640 36660 6680 36720
rect 6740 36660 6780 36720
rect 6840 36660 6880 36720
rect 6940 36660 6980 36720
rect 7040 36660 7080 36720
rect 7140 36660 7180 36720
rect 7240 36660 7280 36720
rect 7340 36660 7380 36720
rect 7440 36660 7480 36720
rect 7540 36660 7580 36720
rect 7640 36660 7680 36720
rect 7740 36660 7780 36720
rect 7840 36660 7880 36720
rect 7940 36660 7980 36720
rect 8040 36660 8080 36720
rect 8140 36660 8180 36720
rect 8240 36660 8280 36720
rect 8340 36660 8380 36720
rect 8440 36660 8480 36720
rect 8540 36660 8580 36720
rect 8640 36660 8680 36720
rect 8740 36660 8780 36720
rect 8840 36660 8880 36720
rect 8940 36660 8980 36720
rect 9040 36660 9080 36720
rect 9140 36660 9180 36720
rect 9240 36660 9280 36720
rect 9340 36660 9380 36720
rect 9440 36660 9480 36720
rect 9540 36660 9580 36720
rect 9640 36660 9680 36720
rect 9740 36660 9780 36720
rect 9840 36660 9880 36720
rect 9940 36660 9980 36720
rect 10040 36660 10080 36720
rect 10140 36660 10180 36720
rect 10240 36660 10280 36720
rect 10340 36660 10380 36720
rect 10440 36660 10480 36720
rect 10540 36660 10580 36720
rect 10640 36660 10680 36720
rect 10740 36660 10780 36720
rect 10840 36660 10930 36720
rect 6340 36650 10930 36660
rect 12920 37200 24910 37260
rect 12920 36400 12970 37200
rect 13760 36400 13970 37200
rect 14760 36400 24910 37200
rect 12920 36340 24910 36400
rect 8660 35470 8780 35500
rect 8660 35460 11690 35470
rect 8660 35370 8680 35460
rect 8760 35370 11690 35460
rect 8660 35360 11690 35370
rect 8660 35330 8780 35360
rect 3670 34990 3840 35010
rect 3670 34940 3760 34990
rect 3810 34940 3840 34990
rect 3670 34920 3840 34940
rect 4530 35000 4650 35010
rect 4530 34930 4560 35000
rect 4620 34930 4650 35000
rect 9050 34950 9110 34970
rect 4530 34920 4650 34930
rect 3670 33630 3730 34920
rect 6190 34910 9060 34950
rect 9100 34910 9110 34950
rect 5300 34870 5530 34890
rect 6190 34870 6260 34910
rect 9050 34890 9110 34910
rect 5300 34820 5310 34870
rect 5360 34820 5420 34870
rect 5470 34820 5530 34870
rect 5300 34800 5530 34820
rect 6120 34860 6260 34870
rect 6710 34860 6770 34870
rect 6120 34810 6190 34860
rect 6240 34850 6410 34860
rect 6240 34810 6340 34850
rect 6380 34810 6410 34850
rect 6120 34800 6410 34810
rect 6520 34850 6770 34860
rect 8790 34850 8850 34860
rect 6520 34810 6640 34850
rect 6680 34810 6720 34850
rect 6760 34810 6770 34850
rect 6520 34800 6770 34810
rect 6710 34790 6770 34800
rect 7070 34840 7370 34850
rect 7070 34800 7220 34840
rect 7260 34800 7300 34840
rect 7340 34800 7370 34840
rect 7070 34790 7370 34800
rect 7480 34840 7750 34850
rect 7480 34800 7600 34840
rect 7640 34800 7680 34840
rect 7720 34800 7750 34840
rect 7480 34790 7750 34800
rect 7860 34840 8130 34850
rect 7860 34800 7980 34840
rect 8020 34800 8060 34840
rect 8100 34800 8130 34840
rect 7860 34790 8130 34800
rect 8240 34840 8510 34850
rect 8240 34800 8360 34840
rect 8400 34800 8440 34840
rect 8480 34800 8510 34840
rect 8240 34790 8510 34800
rect 8620 34840 8850 34850
rect 8620 34800 8690 34840
rect 8730 34800 8800 34840
rect 8840 34800 8850 34840
rect 8620 34790 8850 34800
rect 9150 34840 9450 34850
rect 9150 34800 9300 34840
rect 9340 34800 9380 34840
rect 9420 34800 9450 34840
rect 9150 34790 9450 34800
rect 9560 34840 9830 34850
rect 9560 34800 9680 34840
rect 9720 34800 9760 34840
rect 9800 34800 9830 34840
rect 9560 34790 9830 34800
rect 9940 34840 10210 34850
rect 9940 34800 10060 34840
rect 10100 34800 10140 34840
rect 10180 34800 10210 34840
rect 9940 34790 10210 34800
rect 10320 34840 10590 34850
rect 10320 34800 10440 34840
rect 10480 34800 10520 34840
rect 10560 34800 10590 34840
rect 10320 34790 10590 34800
rect 10700 34840 10880 34850
rect 10700 34800 10820 34840
rect 10860 34800 10880 34840
rect 10700 34790 10880 34800
rect 8790 34780 8850 34790
rect 7170 34190 7230 34210
rect 10820 34190 10860 34790
rect 7170 34150 7180 34190
rect 7220 34150 10860 34190
rect 7170 34130 7230 34150
rect 6270 34040 10880 34050
rect 6270 33980 6380 34040
rect 6440 33980 6480 34040
rect 6540 33980 6580 34040
rect 6640 33980 6680 34040
rect 6740 33980 6780 34040
rect 6840 33980 6880 34040
rect 6940 33980 6980 34040
rect 7040 33980 7080 34040
rect 7140 33980 7180 34040
rect 7240 33980 7280 34040
rect 7340 33980 7380 34040
rect 7440 33980 7480 34040
rect 7540 33980 7580 34040
rect 7640 33980 7680 34040
rect 7740 33980 7780 34040
rect 7840 33980 7880 34040
rect 7940 33980 7980 34040
rect 8040 33980 8080 34040
rect 8140 33980 8180 34040
rect 8240 33980 8280 34040
rect 8340 33980 8380 34040
rect 8440 33980 8480 34040
rect 8540 33980 8580 34040
rect 8640 33980 8680 34040
rect 8740 33980 8780 34040
rect 8840 33980 8880 34040
rect 8940 33980 8980 34040
rect 9040 33980 9080 34040
rect 9140 33980 9180 34040
rect 9240 33980 9280 34040
rect 9340 33980 9380 34040
rect 9440 33980 9480 34040
rect 9540 33980 9580 34040
rect 9640 33980 9680 34040
rect 9740 33980 9780 34040
rect 9840 33980 9880 34040
rect 9940 33980 9980 34040
rect 10040 33980 10080 34040
rect 10140 33980 10180 34040
rect 10240 33980 10280 34040
rect 10340 33980 10380 34040
rect 10440 33980 10480 34040
rect 10540 33980 10580 34040
rect 10640 33980 10680 34040
rect 10740 33980 10780 34040
rect 10840 33980 10880 34040
rect 6270 33970 10880 33980
rect 6270 33630 10920 33970
rect 2070 33620 10920 33630
rect 2070 33560 3810 33620
rect 3870 33560 3910 33620
rect 3970 33560 4010 33620
rect 4070 33560 4110 33620
rect 4170 33560 4210 33620
rect 4270 33560 4310 33620
rect 4370 33560 4410 33620
rect 4470 33560 4510 33620
rect 4570 33560 4610 33620
rect 4670 33560 4710 33620
rect 4770 33560 4810 33620
rect 4870 33560 4910 33620
rect 4970 33560 5010 33620
rect 5070 33560 5110 33620
rect 5170 33560 5210 33620
rect 5270 33560 5310 33620
rect 5370 33560 5410 33620
rect 5470 33560 5510 33620
rect 5570 33560 5610 33620
rect 5670 33560 5710 33620
rect 5770 33560 5810 33620
rect 5870 33560 5910 33620
rect 5970 33560 6010 33620
rect 6070 33560 6110 33620
rect 6170 33560 10920 33620
rect 2070 33360 10920 33560
rect 2070 32670 2120 33360
rect 2950 32670 3150 33360
rect 3980 32670 4180 33360
rect 5010 32670 5210 33360
rect 6040 32670 6240 33360
rect 7070 32670 7270 33360
rect 8100 32670 8300 33360
rect 9130 32670 9330 33360
rect 10870 32670 10920 33360
rect 2070 32620 10920 32670
rect 2070 32480 11240 32540
rect 2070 31790 2120 32480
rect 2950 31790 3150 32480
rect 3980 31790 4180 32480
rect 5010 31790 5210 32480
rect 6040 31790 6240 32480
rect 7070 31790 7270 32480
rect 8100 31790 8300 32480
rect 9130 31790 9330 32480
rect 10160 31790 10360 32480
rect 11190 31790 11240 32480
rect 2070 31740 11240 31790
rect 2170 31730 11240 31740
rect 2170 31670 2210 31730
rect 2270 31670 2310 31730
rect 2370 31670 2410 31730
rect 2470 31670 2510 31730
rect 2570 31670 2610 31730
rect 2670 31670 2710 31730
rect 2770 31670 2810 31730
rect 2870 31670 2910 31730
rect 2970 31670 3010 31730
rect 3070 31670 3110 31730
rect 3170 31670 3210 31730
rect 3270 31670 3310 31730
rect 3370 31670 3410 31730
rect 3470 31670 3510 31730
rect 3570 31670 3610 31730
rect 3670 31670 3710 31730
rect 3770 31670 3810 31730
rect 3870 31670 3910 31730
rect 3970 31670 4010 31730
rect 4070 31670 4110 31730
rect 4170 31670 4210 31730
rect 4270 31670 4310 31730
rect 4370 31670 4410 31730
rect 4470 31670 4510 31730
rect 4570 31670 4610 31730
rect 4670 31670 4710 31730
rect 4770 31670 4810 31730
rect 4870 31670 4910 31730
rect 4970 31670 5010 31730
rect 5070 31670 5110 31730
rect 5170 31670 5210 31730
rect 5270 31670 5310 31730
rect 5370 31670 5410 31730
rect 5470 31670 5510 31730
rect 5570 31670 5610 31730
rect 5670 31670 5710 31730
rect 5770 31670 5810 31730
rect 5870 31670 5910 31730
rect 5970 31670 6010 31730
rect 6070 31670 6110 31730
rect 6170 31670 6210 31730
rect 6270 31670 11240 31730
rect 2170 31660 11240 31670
rect 6380 31380 11240 31660
rect 6380 31320 6470 31380
rect 6530 31320 6580 31380
rect 6640 31320 6690 31380
rect 6750 31320 6800 31380
rect 6860 31320 6910 31380
rect 6970 31320 7020 31380
rect 7080 31320 7130 31380
rect 7190 31320 7240 31380
rect 7300 31320 7350 31380
rect 7410 31320 7460 31380
rect 7520 31320 7570 31380
rect 7630 31320 7680 31380
rect 7740 31320 7790 31380
rect 7850 31320 7900 31380
rect 7960 31320 8010 31380
rect 8070 31320 8120 31380
rect 8180 31320 8230 31380
rect 8290 31320 8340 31380
rect 8400 31320 8450 31380
rect 8510 31320 8560 31380
rect 8620 31320 8670 31380
rect 8730 31320 8780 31380
rect 8840 31320 8890 31380
rect 8950 31320 9000 31380
rect 9060 31320 9110 31380
rect 9170 31320 9220 31380
rect 9280 31320 9330 31380
rect 9390 31320 9440 31380
rect 9500 31320 9550 31380
rect 9610 31320 9660 31380
rect 9720 31320 9770 31380
rect 9830 31320 9880 31380
rect 9940 31320 9990 31380
rect 10050 31320 10100 31380
rect 10160 31320 10210 31380
rect 10270 31320 10320 31380
rect 10380 31320 10430 31380
rect 10490 31320 10540 31380
rect 10600 31320 10650 31380
rect 10710 31320 10760 31380
rect 10820 31320 10880 31380
rect 10940 31320 10990 31380
rect 11050 31320 11100 31380
rect 11160 31320 11240 31380
rect 6380 31300 11240 31320
rect 9110 30800 9170 30820
rect 6310 30760 9120 30800
rect 9160 30760 9170 30800
rect 2070 30740 2240 30760
rect 2070 30690 2160 30740
rect 2210 30690 2240 30740
rect 2070 30670 2240 30690
rect 2930 30740 3050 30760
rect 2930 30680 2960 30740
rect 3020 30680 3050 30740
rect 6310 30720 6380 30760
rect 9110 30740 9170 30760
rect 11170 30720 11470 30740
rect 2930 30670 3050 30680
rect 6240 30710 6380 30720
rect 6770 30710 6830 30720
rect 2070 29380 2130 30670
rect 6240 30660 6310 30710
rect 6360 30700 6470 30710
rect 6360 30660 6400 30700
rect 6440 30660 6470 30700
rect 6240 30650 6470 30660
rect 6580 30700 6830 30710
rect 8850 30700 8910 30710
rect 6580 30660 6700 30700
rect 6740 30660 6780 30700
rect 6820 30660 6830 30700
rect 6580 30650 6830 30660
rect 6770 30640 6830 30650
rect 7130 30690 7430 30700
rect 7130 30650 7280 30690
rect 7320 30650 7360 30690
rect 7400 30650 7430 30690
rect 7130 30640 7430 30650
rect 7540 30690 7810 30700
rect 7540 30650 7660 30690
rect 7700 30650 7740 30690
rect 7780 30650 7810 30690
rect 7540 30640 7810 30650
rect 7920 30690 8190 30700
rect 7920 30650 8040 30690
rect 8080 30650 8120 30690
rect 8160 30650 8190 30690
rect 7920 30640 8190 30650
rect 8300 30690 8570 30700
rect 8300 30650 8420 30690
rect 8460 30650 8500 30690
rect 8540 30650 8570 30690
rect 8300 30640 8570 30650
rect 8680 30690 8910 30700
rect 8680 30650 8750 30690
rect 8790 30650 8860 30690
rect 8900 30650 8910 30690
rect 8680 30640 8910 30650
rect 9210 30690 9510 30700
rect 9210 30650 9360 30690
rect 9400 30650 9440 30690
rect 9480 30650 9510 30690
rect 9210 30640 9510 30650
rect 9620 30690 9890 30700
rect 9620 30650 9740 30690
rect 9780 30650 9820 30690
rect 9860 30650 9890 30690
rect 9620 30640 9890 30650
rect 10000 30690 10270 30700
rect 10000 30650 10120 30690
rect 10160 30650 10200 30690
rect 10240 30650 10270 30690
rect 10000 30640 10270 30650
rect 10380 30690 10650 30700
rect 10380 30650 10500 30690
rect 10540 30650 10580 30690
rect 10620 30650 10650 30690
rect 10380 30640 10650 30650
rect 10760 30690 11030 30700
rect 10760 30650 10880 30690
rect 10920 30650 10960 30690
rect 11000 30650 11030 30690
rect 10760 30640 11030 30650
rect 11170 30660 11240 30720
rect 11300 30660 11470 30720
rect 11170 30640 11470 30660
rect 8850 30630 8910 30640
rect 3700 30610 3800 30620
rect 4520 30610 4790 30620
rect 3700 30600 3930 30610
rect 3700 30560 3730 30600
rect 3770 30560 3820 30600
rect 3860 30560 3930 30600
rect 3700 30550 3930 30560
rect 4520 30560 4590 30610
rect 4640 30560 4680 30610
rect 4730 30560 4790 30610
rect 4520 30550 4790 30560
rect 5380 30610 5650 30620
rect 5380 30560 5450 30610
rect 5500 30560 5540 30610
rect 5590 30560 5650 30610
rect 5380 30550 5650 30560
rect 3700 30540 3800 30550
rect 7230 30040 7290 30060
rect 10880 30040 10920 30640
rect 7230 30000 7240 30040
rect 7280 30000 10920 30040
rect 7230 29980 7290 30000
rect 6330 29900 11240 29910
rect 6330 29840 6440 29900
rect 6500 29840 6540 29900
rect 6600 29840 6640 29900
rect 6700 29840 6740 29900
rect 6800 29840 6840 29900
rect 6900 29840 6940 29900
rect 7000 29840 7040 29900
rect 7100 29840 7140 29900
rect 7200 29840 7240 29900
rect 7300 29840 7340 29900
rect 7400 29840 7440 29900
rect 7500 29840 7540 29900
rect 7600 29840 7640 29900
rect 7700 29840 7740 29900
rect 7800 29840 7840 29900
rect 7900 29840 7940 29900
rect 8000 29840 8040 29900
rect 8100 29840 8140 29900
rect 8200 29840 8240 29900
rect 8300 29840 8340 29900
rect 8400 29840 8440 29900
rect 8500 29840 8540 29900
rect 8600 29840 8640 29900
rect 8700 29840 8740 29900
rect 8800 29840 8840 29900
rect 8900 29840 8940 29900
rect 9000 29840 9040 29900
rect 9100 29840 9140 29900
rect 9200 29840 9240 29900
rect 9300 29840 9340 29900
rect 9400 29840 9440 29900
rect 9500 29840 9540 29900
rect 9600 29840 9640 29900
rect 9700 29840 9740 29900
rect 9800 29840 9840 29900
rect 9900 29840 9940 29900
rect 10000 29840 10040 29900
rect 10100 29840 10140 29900
rect 10200 29840 10240 29900
rect 10300 29840 10340 29900
rect 10400 29840 10440 29900
rect 10500 29840 10540 29900
rect 10600 29840 10640 29900
rect 10700 29840 10740 29900
rect 10800 29840 10840 29900
rect 10900 29840 10940 29900
rect 11000 29840 11040 29900
rect 11100 29840 11140 29900
rect 11200 29840 11240 29900
rect 6330 29380 11240 29840
rect 2070 29370 11240 29380
rect 2070 29310 2210 29370
rect 2270 29310 2310 29370
rect 2370 29310 2410 29370
rect 2470 29310 2510 29370
rect 2570 29310 2610 29370
rect 2670 29310 2710 29370
rect 2770 29310 2810 29370
rect 2870 29310 2910 29370
rect 2970 29310 3010 29370
rect 3070 29310 3110 29370
rect 3170 29310 3210 29370
rect 3270 29310 3310 29370
rect 3370 29310 3410 29370
rect 3470 29310 3510 29370
rect 3570 29310 3610 29370
rect 3670 29310 3710 29370
rect 3770 29310 3810 29370
rect 3870 29310 3910 29370
rect 3970 29310 4010 29370
rect 4070 29310 4110 29370
rect 4170 29310 4210 29370
rect 4270 29310 4310 29370
rect 4370 29310 4410 29370
rect 4470 29310 4510 29370
rect 4570 29310 4610 29370
rect 4670 29310 4710 29370
rect 4770 29310 4810 29370
rect 4870 29310 4910 29370
rect 4970 29310 5010 29370
rect 5070 29310 5110 29370
rect 5170 29310 5210 29370
rect 5270 29310 5310 29370
rect 5370 29310 5410 29370
rect 5470 29310 5510 29370
rect 5570 29310 5610 29370
rect 5670 29310 5710 29370
rect 5770 29310 5810 29370
rect 5870 29310 5910 29370
rect 5970 29310 6010 29370
rect 6070 29310 6110 29370
rect 6170 29310 6210 29370
rect 6270 29310 11240 29370
rect 2070 29000 11240 29310
rect 2070 28310 2120 29000
rect 2950 28310 3150 29000
rect 3980 28310 4180 29000
rect 5010 28310 5210 29000
rect 6040 28310 6240 29000
rect 7070 28310 7270 29000
rect 8100 28310 8300 29000
rect 9130 28310 9330 29000
rect 10160 28310 10360 29000
rect 11190 28310 11240 29000
rect 2070 28260 11240 28310
rect 5360 28100 5500 28120
rect 5360 27990 5380 28100
rect 5480 27990 5500 28100
rect 11370 28030 11470 30640
rect 5360 27970 5500 27990
rect 5380 10420 5480 27970
rect 6740 27940 11470 28030
rect 5590 27820 5730 27840
rect 5590 27710 5610 27820
rect 5710 27710 5730 27820
rect 5590 27690 5730 27710
rect 5610 12730 5710 27690
rect 6280 25560 6380 25580
rect 6280 25500 6300 25560
rect 6360 25500 6380 25560
rect 6280 25480 6380 25500
rect 6740 25210 6820 27940
rect 11570 27910 11690 35360
rect 12920 33100 13830 36340
rect 15180 36270 15220 36340
rect 15280 36270 15320 36340
rect 15380 36270 15420 36340
rect 15480 36270 15520 36340
rect 15580 36270 15620 36340
rect 15680 36270 15720 36340
rect 15780 36270 15820 36340
rect 15880 36270 15920 36340
rect 15980 36270 16020 36340
rect 16080 36270 16120 36340
rect 16180 36270 16220 36340
rect 16280 36270 16320 36340
rect 16380 36270 16420 36340
rect 16480 36270 16520 36340
rect 16580 36270 16620 36340
rect 16680 36270 16720 36340
rect 16780 36270 16820 36340
rect 16880 36270 16920 36340
rect 16980 36270 17020 36340
rect 17080 36270 17120 36340
rect 17180 36270 17220 36340
rect 17280 36270 17320 36340
rect 17380 36270 17420 36340
rect 17480 36270 17520 36340
rect 17580 36270 17620 36340
rect 17680 36270 17720 36340
rect 17780 36270 17820 36340
rect 17880 36270 17920 36340
rect 17980 36270 18020 36340
rect 18080 36270 18120 36340
rect 18180 36270 18220 36340
rect 18280 36270 18320 36340
rect 18380 36270 18420 36340
rect 18480 36270 18520 36340
rect 18580 36270 18620 36340
rect 18680 36270 18720 36340
rect 18780 36270 18820 36340
rect 18880 36270 18920 36340
rect 18980 36270 19020 36340
rect 19080 36270 19120 36340
rect 19180 36270 19220 36340
rect 19280 36270 19320 36340
rect 19380 36270 19420 36340
rect 19480 36270 19520 36340
rect 19580 36270 19620 36340
rect 19680 36270 19720 36340
rect 19780 36270 19820 36340
rect 19880 36270 19920 36340
rect 19980 36270 20020 36340
rect 20080 36270 20120 36340
rect 20180 36270 20220 36340
rect 20280 36270 20320 36340
rect 20380 36270 20420 36340
rect 20480 36270 20520 36340
rect 20580 36270 20620 36340
rect 20680 36270 20720 36340
rect 20780 36270 20820 36340
rect 20880 36270 20920 36340
rect 20980 36270 21020 36340
rect 21080 36270 21120 36340
rect 21180 36270 21220 36340
rect 21280 36270 21320 36340
rect 21380 36270 21420 36340
rect 21480 36270 21520 36340
rect 21580 36270 21620 36340
rect 21680 36270 21720 36340
rect 21780 36270 21820 36340
rect 21880 36270 21920 36340
rect 21980 36270 22020 36340
rect 22080 36270 22120 36340
rect 22180 36270 22220 36340
rect 22280 36270 22320 36340
rect 22380 36270 22420 36340
rect 22480 36270 22520 36340
rect 22580 36270 22620 36340
rect 22680 36270 22720 36340
rect 22780 36270 22820 36340
rect 22880 36270 22920 36340
rect 22980 36270 23020 36340
rect 23080 36270 23120 36340
rect 23180 36270 23220 36340
rect 23280 36270 23320 36340
rect 23380 36270 23420 36340
rect 23480 36270 23520 36340
rect 23580 36270 23620 36340
rect 23680 36270 23720 36340
rect 23780 36270 23820 36340
rect 23880 36270 23920 36340
rect 23980 36270 24020 36340
rect 24080 36270 24120 36340
rect 24180 36270 24220 36340
rect 24280 36270 24320 36340
rect 24380 36270 24420 36340
rect 24480 36270 24520 36340
rect 24580 36270 24620 36340
rect 24680 36270 24720 36340
rect 24780 36270 24820 36340
rect 24880 36270 24910 36340
rect 15180 36260 24910 36270
rect 15220 36120 15280 36260
rect 17220 36150 18350 36200
rect 15160 36110 15340 36120
rect 15160 36050 15200 36110
rect 15300 36050 15340 36110
rect 15440 36110 15520 36120
rect 15440 36070 15460 36110
rect 15500 36070 15520 36110
rect 15440 36060 15520 36070
rect 17220 36060 17300 36150
rect 15160 36040 15340 36050
rect 15860 35980 17300 36060
rect 15860 35880 15910 35980
rect 15860 35830 16010 35880
rect 15550 35630 15660 35640
rect 15550 35570 15570 35630
rect 15640 35570 15660 35630
rect 15550 35560 15660 35570
rect 15760 35630 15930 35640
rect 15760 35570 15790 35630
rect 15900 35570 15930 35630
rect 15760 35560 15930 35570
rect 15450 35520 15510 35540
rect 15960 35520 16010 35830
rect 15450 35480 15460 35520
rect 15500 35480 16010 35520
rect 16430 35490 16530 35510
rect 15450 35460 15510 35480
rect 16430 35430 16450 35490
rect 16510 35430 16530 35490
rect 17120 35490 17200 35500
rect 17560 35490 17780 35500
rect 17120 35450 17140 35490
rect 17180 35450 17300 35490
rect 17120 35440 17200 35450
rect 16430 35410 16530 35430
rect 17250 35330 17300 35450
rect 17560 35450 17580 35490
rect 17620 35450 17720 35490
rect 17760 35450 17780 35490
rect 17560 35440 17780 35450
rect 18020 35490 18100 35500
rect 18020 35450 18040 35490
rect 18080 35450 18100 35490
rect 18020 35440 18100 35450
rect 17640 35360 17700 35440
rect 17220 35310 17330 35330
rect 17220 35240 17240 35310
rect 17310 35240 17330 35310
rect 17640 35320 17650 35360
rect 17690 35320 17700 35360
rect 18260 35320 18350 36150
rect 20710 36170 20810 36190
rect 20710 36090 20730 36170
rect 20790 36090 20810 36170
rect 20710 36070 20810 36090
rect 20740 35930 20780 36070
rect 20710 35910 20810 35930
rect 20710 35830 20730 35910
rect 20790 35830 20810 35910
rect 20710 35810 20810 35830
rect 19870 35520 20080 35530
rect 18500 35490 18720 35500
rect 18500 35450 18520 35490
rect 18560 35450 18660 35490
rect 18700 35450 18720 35490
rect 18500 35440 18720 35450
rect 18960 35490 19040 35500
rect 19750 35490 19830 35500
rect 18960 35450 18980 35490
rect 19020 35450 19040 35490
rect 18960 35440 19040 35450
rect 19580 35450 19770 35490
rect 19810 35450 19830 35490
rect 19870 35480 20020 35520
rect 20060 35480 20080 35520
rect 24830 35520 25040 35530
rect 19870 35470 20080 35480
rect 21330 35490 21490 35500
rect 17640 35300 17700 35320
rect 18220 35300 18350 35320
rect 18580 35360 18640 35440
rect 18580 35320 18590 35360
rect 18630 35320 18640 35360
rect 18580 35300 18640 35320
rect 17220 35220 17330 35240
rect 18220 35230 18270 35300
rect 18340 35280 18350 35300
rect 18340 35270 18360 35280
rect 18340 35230 18620 35270
rect 17250 34610 17300 35220
rect 18220 35210 18350 35230
rect 17850 35200 18270 35210
rect 17850 35160 17870 35200
rect 17910 35160 18270 35200
rect 17850 35150 18270 35160
rect 17450 34900 17530 34910
rect 17450 34860 17470 34900
rect 17510 34860 17530 34900
rect 17450 34850 17530 34860
rect 18390 34900 18470 34910
rect 18390 34860 18410 34900
rect 18450 34860 18470 34900
rect 18570 34900 18620 35230
rect 19580 34970 19640 35450
rect 19750 35440 19830 35450
rect 21330 35450 21430 35490
rect 21470 35450 21490 35490
rect 21330 35440 21490 35450
rect 22080 35490 22160 35500
rect 22520 35490 22740 35500
rect 22080 35450 22100 35490
rect 22140 35450 22250 35490
rect 22080 35440 22160 35450
rect 20120 35370 20620 35390
rect 20120 35330 20210 35370
rect 20250 35330 20620 35370
rect 20120 35310 20620 35330
rect 18970 34950 19200 34970
rect 19310 34950 19370 34970
rect 18970 34910 19130 34950
rect 19170 34910 19320 34950
rect 19360 34910 19370 34950
rect 18680 34900 18760 34910
rect 18570 34860 18700 34900
rect 18740 34860 18760 34900
rect 18970 34890 19200 34910
rect 19310 34890 19370 34910
rect 19410 34950 19640 34970
rect 19410 34910 19520 34950
rect 19560 34910 19640 34950
rect 19410 34890 19640 34910
rect 18390 34850 18470 34860
rect 18680 34850 18760 34860
rect 17470 34820 17510 34850
rect 18410 34820 18450 34850
rect 17470 34780 18450 34820
rect 17470 34610 17510 34780
rect 17250 34560 17510 34610
rect 17860 34670 18860 34710
rect 17860 34370 17920 34670
rect 18290 34620 18390 34670
rect 18290 34540 18310 34620
rect 18370 34540 18390 34620
rect 18290 34530 18390 34540
rect 18800 34370 18860 34670
rect 19580 34660 19640 34890
rect 19730 34810 19830 34830
rect 19730 34750 19750 34810
rect 19810 34750 19830 34810
rect 19870 34820 19930 34830
rect 19870 34810 20080 34820
rect 19870 34770 19880 34810
rect 19920 34770 20020 34810
rect 20060 34770 20080 34810
rect 19870 34760 20080 34770
rect 19870 34750 19930 34760
rect 19730 34730 19830 34750
rect 19750 34660 19830 34670
rect 19580 34620 19770 34660
rect 19810 34620 19830 34660
rect 19580 34450 19640 34620
rect 19750 34610 19830 34620
rect 20540 34530 20620 35310
rect 20900 34960 21000 34980
rect 20900 34900 20920 34960
rect 20980 34900 21000 34960
rect 20900 34880 21000 34900
rect 21140 34950 21240 34970
rect 21330 34950 21370 35440
rect 22210 35330 22250 35450
rect 22520 35450 22540 35490
rect 22580 35450 22680 35490
rect 22720 35450 22740 35490
rect 22520 35440 22740 35450
rect 22980 35490 23060 35500
rect 22980 35450 23000 35490
rect 23040 35450 23060 35490
rect 22980 35440 23060 35450
rect 23460 35490 23680 35500
rect 23460 35450 23480 35490
rect 23520 35450 23620 35490
rect 23660 35450 23680 35490
rect 23460 35440 23680 35450
rect 23920 35490 24000 35500
rect 24710 35490 24790 35500
rect 23920 35450 23940 35490
rect 23980 35450 24000 35490
rect 23920 35440 24000 35450
rect 24550 35450 24730 35490
rect 24770 35450 24790 35490
rect 24830 35480 24980 35520
rect 25020 35480 25040 35520
rect 24830 35470 25040 35480
rect 22600 35360 22660 35440
rect 22180 35310 22290 35330
rect 22180 35240 22200 35310
rect 22270 35240 22290 35310
rect 22600 35320 22610 35360
rect 22650 35320 22660 35360
rect 22600 35300 22660 35320
rect 23540 35360 23600 35440
rect 23540 35320 23550 35360
rect 23590 35320 23600 35360
rect 23540 35300 23600 35320
rect 22180 35220 22290 35240
rect 23180 35240 23600 35270
rect 21140 34910 21190 34950
rect 21230 34910 21370 34950
rect 21140 34890 21240 34910
rect 22210 34690 22250 35220
rect 23180 35210 23520 35240
rect 22810 35200 22890 35210
rect 23180 35200 23230 35210
rect 22810 35160 22830 35200
rect 22870 35160 23230 35200
rect 23510 35170 23520 35210
rect 23590 35170 23600 35240
rect 22810 35150 22890 35160
rect 23510 35150 23600 35170
rect 22410 34900 22490 34910
rect 22410 34860 22430 34900
rect 22470 34860 22490 34900
rect 22410 34850 22490 34860
rect 23350 34900 23430 34910
rect 23350 34860 23370 34900
rect 23410 34860 23430 34900
rect 23530 34900 23580 35150
rect 24550 34970 24600 35450
rect 24710 35440 24790 35450
rect 25080 35370 26430 35390
rect 25080 35330 25170 35370
rect 25210 35330 26430 35370
rect 25080 35310 26430 35330
rect 23930 34950 24160 34970
rect 24270 34950 24330 34970
rect 23930 34910 24090 34950
rect 24130 34910 24280 34950
rect 24320 34910 24330 34950
rect 23640 34900 23720 34910
rect 23530 34860 23660 34900
rect 23700 34860 23720 34900
rect 23930 34890 24160 34910
rect 24270 34890 24330 34910
rect 24370 34950 24600 34970
rect 24370 34910 24480 34950
rect 24520 34910 24600 34950
rect 24370 34890 24600 34910
rect 23350 34850 23430 34860
rect 23640 34850 23720 34860
rect 22430 34820 22470 34850
rect 23370 34820 23410 34850
rect 22430 34780 23410 34820
rect 22430 34690 22470 34780
rect 22210 34650 22470 34690
rect 22820 34690 23820 34730
rect 20740 34530 20840 34550
rect 20540 34450 20760 34530
rect 20820 34450 20840 34530
rect 19560 34430 19660 34450
rect 20740 34430 20840 34450
rect 17670 34360 18100 34370
rect 17670 34320 17690 34360
rect 17730 34320 17870 34360
rect 17910 34320 18040 34360
rect 18080 34320 18100 34360
rect 17670 34310 18100 34320
rect 18610 34360 19040 34370
rect 18610 34320 18630 34360
rect 18670 34320 18810 34360
rect 18850 34320 18980 34360
rect 19020 34320 19040 34360
rect 19560 34350 19580 34430
rect 19640 34350 19660 34430
rect 22820 34370 22880 34690
rect 23220 34550 23320 34690
rect 23220 34470 23240 34550
rect 23300 34470 23320 34550
rect 23220 34460 23320 34470
rect 23760 34370 23820 34690
rect 24550 34660 24600 34890
rect 24690 34810 24790 34830
rect 24690 34750 24710 34810
rect 24770 34750 24790 34810
rect 24830 34820 24890 34830
rect 24830 34810 25040 34820
rect 24830 34770 24840 34810
rect 24880 34770 24980 34810
rect 25020 34770 25040 34810
rect 24830 34760 25040 34770
rect 24830 34750 24890 34760
rect 24690 34730 24790 34750
rect 24710 34660 24790 34670
rect 24550 34620 24730 34660
rect 24770 34620 24790 34660
rect 19560 34330 19660 34350
rect 22630 34360 23060 34370
rect 18610 34310 19040 34320
rect 22630 34320 22650 34360
rect 22690 34320 22830 34360
rect 22870 34320 23000 34360
rect 23040 34320 23060 34360
rect 22630 34310 23060 34320
rect 23570 34360 24000 34370
rect 23570 34320 23590 34360
rect 23630 34320 23770 34360
rect 23810 34320 23940 34360
rect 23980 34320 24000 34360
rect 23570 34310 24000 34320
rect 24550 34330 24600 34620
rect 24710 34610 24790 34620
rect 24930 34380 25030 34400
rect 24930 34330 24950 34380
rect 24550 34300 24950 34330
rect 25010 34300 25030 34380
rect 24550 34280 25030 34300
rect 16460 34200 25450 34210
rect 16460 34130 16510 34200
rect 16570 34130 16610 34200
rect 16670 34130 16710 34200
rect 16770 34130 16810 34200
rect 16870 34130 16910 34200
rect 16970 34130 17010 34200
rect 17070 34130 17110 34200
rect 17170 34130 17210 34200
rect 17270 34130 17310 34200
rect 17370 34130 17410 34200
rect 17470 34130 17510 34200
rect 17570 34130 17610 34200
rect 17670 34130 17710 34200
rect 17770 34130 17810 34200
rect 17870 34130 17910 34200
rect 17970 34130 18010 34200
rect 18070 34130 18110 34200
rect 18170 34130 18210 34200
rect 18270 34130 18310 34200
rect 18370 34130 18410 34200
rect 18470 34130 18510 34200
rect 18570 34130 18610 34200
rect 18670 34130 18710 34200
rect 18770 34130 18810 34200
rect 18870 34130 18910 34200
rect 18970 34130 19010 34200
rect 19070 34130 19110 34200
rect 19170 34130 19210 34200
rect 19270 34130 19310 34200
rect 19370 34130 19410 34200
rect 19470 34130 19510 34200
rect 19570 34130 19610 34200
rect 19670 34130 19710 34200
rect 19770 34130 19810 34200
rect 19870 34130 19910 34200
rect 19970 34130 20010 34200
rect 20070 34130 20110 34200
rect 20170 34130 20210 34200
rect 20270 34130 20310 34200
rect 20370 34130 20410 34200
rect 20470 34130 20510 34200
rect 20570 34130 20610 34200
rect 20670 34130 20710 34200
rect 20770 34130 20810 34200
rect 20870 34130 20910 34200
rect 20970 34130 21010 34200
rect 21070 34130 21110 34200
rect 21170 34130 21210 34200
rect 21270 34130 21310 34200
rect 21370 34130 21410 34200
rect 21470 34130 21510 34200
rect 21570 34130 21610 34200
rect 21670 34130 21710 34200
rect 21770 34130 21810 34200
rect 21870 34130 21910 34200
rect 21970 34130 22010 34200
rect 22070 34130 22110 34200
rect 22170 34130 22210 34200
rect 22270 34130 22310 34200
rect 22370 34130 22410 34200
rect 22470 34130 22510 34200
rect 22570 34130 22610 34200
rect 22670 34130 22710 34200
rect 22770 34130 22810 34200
rect 22870 34130 22910 34200
rect 22970 34130 23010 34200
rect 23070 34130 23110 34200
rect 23170 34130 23210 34200
rect 23270 34130 23310 34200
rect 23370 34130 23410 34200
rect 23470 34130 23510 34200
rect 23570 34130 23620 34200
rect 23680 34130 23720 34200
rect 23780 34130 23820 34200
rect 23880 34130 23920 34200
rect 23980 34130 24020 34200
rect 24080 34130 24120 34200
rect 24180 34130 24220 34200
rect 24280 34130 24320 34200
rect 24380 34130 24420 34200
rect 24480 34130 24520 34200
rect 24580 34130 24620 34200
rect 24680 34130 24720 34200
rect 24780 34130 24820 34200
rect 24880 34130 24920 34200
rect 24980 34130 25020 34200
rect 25080 34130 25120 34200
rect 25180 34130 25220 34200
rect 25280 34130 25320 34200
rect 25380 34130 25450 34200
rect 16460 34120 25450 34130
rect 15100 34060 25450 34120
rect 15100 33250 22440 34060
rect 23080 33250 25450 34060
rect 15100 33190 25450 33250
rect 12920 32480 25450 33100
rect 13728 32460 13888 32480
rect 13728 32420 13768 32460
rect 13848 32420 13888 32460
rect 13728 32400 13888 32420
rect 14098 32380 14178 32390
rect 14098 32340 14118 32380
rect 14158 32340 14178 32380
rect 14098 32330 14178 32340
rect 15630 32310 15730 32340
rect 14680 32250 15650 32310
rect 15710 32250 15730 32310
rect 14370 32010 14540 32020
rect 14370 31950 14400 32010
rect 14510 31950 14540 32010
rect 13988 31940 14068 31950
rect 14370 31940 14540 31950
rect 13988 31900 14008 31940
rect 14048 31900 14068 31940
rect 13988 31890 14068 31900
rect 14208 31890 14288 31900
rect 14438 31890 14478 31940
rect 14208 31850 14228 31890
rect 14268 31850 14478 31890
rect 14208 31840 14288 31850
rect 14108 31790 14168 31810
rect 14680 31790 14730 32250
rect 15630 32220 15730 32250
rect 16030 32190 25450 32480
rect 16030 32180 25410 32190
rect 16030 32110 16120 32180
rect 16180 32110 16220 32180
rect 16280 32110 16320 32180
rect 16380 32110 16420 32180
rect 16480 32110 16520 32180
rect 16580 32110 16620 32180
rect 16680 32110 16720 32180
rect 16780 32110 16820 32180
rect 16880 32110 16920 32180
rect 16980 32110 17020 32180
rect 17080 32110 17120 32180
rect 17180 32110 17220 32180
rect 17280 32110 17320 32180
rect 17380 32110 17420 32180
rect 17480 32110 17520 32180
rect 17580 32110 17620 32180
rect 17680 32110 17720 32180
rect 17780 32110 17820 32180
rect 17880 32110 17920 32180
rect 17980 32110 18020 32180
rect 18080 32110 18120 32180
rect 18180 32110 18220 32180
rect 18280 32110 18320 32180
rect 18380 32110 18420 32180
rect 18480 32110 18520 32180
rect 18580 32110 18620 32180
rect 18680 32110 18720 32180
rect 18780 32110 18820 32180
rect 18880 32110 18920 32180
rect 18980 32110 19020 32180
rect 19080 32110 19120 32180
rect 19180 32110 19220 32180
rect 19280 32110 19320 32180
rect 19380 32110 19420 32180
rect 19480 32110 19520 32180
rect 19580 32110 19620 32180
rect 19680 32110 19720 32180
rect 19780 32110 19820 32180
rect 19880 32110 19920 32180
rect 19980 32110 20020 32180
rect 20080 32110 20120 32180
rect 20180 32110 20220 32180
rect 20280 32110 20320 32180
rect 20380 32110 20420 32180
rect 20480 32110 20520 32180
rect 20580 32110 20620 32180
rect 20680 32110 20720 32180
rect 20780 32110 20820 32180
rect 20880 32110 20920 32180
rect 20980 32110 21020 32180
rect 21080 32110 21120 32180
rect 21180 32110 21220 32180
rect 21280 32110 21320 32180
rect 21380 32110 21420 32180
rect 21480 32110 21520 32180
rect 21580 32110 21620 32180
rect 21680 32110 21720 32180
rect 21780 32110 21820 32180
rect 21880 32110 21920 32180
rect 21980 32110 22020 32180
rect 22080 32110 22120 32180
rect 22180 32110 22220 32180
rect 22280 32110 22320 32180
rect 22380 32110 22420 32180
rect 22480 32110 22520 32180
rect 22580 32110 22620 32180
rect 22680 32110 22720 32180
rect 22780 32110 22820 32180
rect 22880 32110 22920 32180
rect 22980 32110 23020 32180
rect 23080 32110 23120 32180
rect 23180 32110 23220 32180
rect 23280 32110 23320 32180
rect 23380 32110 23420 32180
rect 23480 32110 23520 32180
rect 23580 32110 23620 32180
rect 23680 32110 23720 32180
rect 23780 32110 23820 32180
rect 23880 32110 23920 32180
rect 23980 32110 24020 32180
rect 24080 32110 24120 32180
rect 24180 32110 24220 32180
rect 24280 32110 24320 32180
rect 24380 32110 24420 32180
rect 24480 32110 24520 32180
rect 24580 32110 24620 32180
rect 24680 32110 24720 32180
rect 24780 32110 24820 32180
rect 24880 32110 24920 32180
rect 24980 32110 25020 32180
rect 25080 32110 25120 32180
rect 25180 32110 25220 32180
rect 25280 32110 25320 32180
rect 25380 32110 25410 32180
rect 16030 32100 25410 32110
rect 15570 32020 15670 32040
rect 15570 31940 15590 32020
rect 15650 31940 15810 32020
rect 15570 31920 15670 31940
rect 14028 31750 14118 31790
rect 14158 31750 14730 31790
rect 14028 31310 14068 31750
rect 14108 31730 14168 31750
rect 14098 31310 14178 31320
rect 14028 31270 14118 31310
rect 14158 31270 14178 31310
rect 14098 31260 14178 31270
rect 15380 30280 15490 30300
rect 15380 30210 15400 30280
rect 15470 30210 15490 30280
rect 15380 30140 15490 30210
rect 15730 30140 15810 31940
rect 16430 31450 16530 31470
rect 25090 31450 25300 31460
rect 16430 31390 16450 31450
rect 16510 31390 16530 31450
rect 20130 31440 20340 31450
rect 16430 31370 16530 31390
rect 17120 31430 17200 31440
rect 17560 31430 17780 31440
rect 17120 31390 17140 31430
rect 17180 31390 17300 31430
rect 17120 31380 17200 31390
rect 17250 31320 17300 31390
rect 17560 31390 17580 31430
rect 17620 31390 17720 31430
rect 17760 31390 17780 31430
rect 17560 31380 17780 31390
rect 18020 31430 18100 31440
rect 18020 31390 18040 31430
rect 18080 31390 18100 31430
rect 18020 31380 18100 31390
rect 18500 31430 18720 31440
rect 18500 31390 18520 31430
rect 18560 31390 18660 31430
rect 18700 31390 18720 31430
rect 18500 31380 18720 31390
rect 18960 31430 19040 31440
rect 20010 31430 20090 31440
rect 18960 31390 18980 31430
rect 19020 31390 19040 31430
rect 18960 31380 19040 31390
rect 19850 31390 20030 31430
rect 20070 31390 20090 31430
rect 20130 31400 20280 31440
rect 20320 31400 20340 31440
rect 21470 31420 21550 31430
rect 20130 31390 20340 31400
rect 17220 31300 17330 31320
rect 17220 31230 17240 31300
rect 17310 31230 17330 31300
rect 17640 31300 17700 31380
rect 17640 31260 17650 31300
rect 17690 31260 17700 31300
rect 17640 31240 17700 31260
rect 18580 31300 18640 31380
rect 18580 31260 18590 31300
rect 18630 31260 18640 31300
rect 18580 31240 18640 31260
rect 17220 31210 17330 31230
rect 17250 30640 17300 31210
rect 18240 31170 18620 31210
rect 17850 31140 17930 31150
rect 18240 31140 18280 31170
rect 17850 31100 17870 31140
rect 17910 31100 18280 31140
rect 18530 31150 18620 31170
rect 17850 31090 17930 31100
rect 18530 31080 18540 31150
rect 18610 31080 18620 31150
rect 18530 31060 18620 31080
rect 17450 30840 17530 30850
rect 17450 30800 17470 30840
rect 17510 30800 17530 30840
rect 17450 30790 17530 30800
rect 18390 30840 18470 30850
rect 18390 30800 18410 30840
rect 18450 30800 18470 30840
rect 18570 30840 18620 31060
rect 19850 30910 19900 31390
rect 20010 31380 20090 31390
rect 21390 31380 21490 31420
rect 21530 31380 21550 31420
rect 20380 31240 20620 31260
rect 20380 31200 20470 31240
rect 20510 31200 20620 31240
rect 20380 31180 20620 31200
rect 18970 30890 19200 30910
rect 19310 30890 19370 30910
rect 18970 30850 19130 30890
rect 19170 30850 19320 30890
rect 19360 30850 19370 30890
rect 18680 30840 18760 30850
rect 18570 30800 18700 30840
rect 18740 30800 18760 30840
rect 18970 30830 19200 30850
rect 19310 30830 19370 30850
rect 19410 30890 19520 30910
rect 19570 30890 19630 30910
rect 19410 30850 19460 30890
rect 19500 30850 19580 30890
rect 19620 30850 19630 30890
rect 19410 30830 19520 30850
rect 19570 30830 19630 30850
rect 19670 30890 19900 30910
rect 19670 30850 19780 30890
rect 19820 30850 19900 30890
rect 19670 30830 19900 30850
rect 18390 30790 18470 30800
rect 18680 30790 18760 30800
rect 17470 30760 17510 30790
rect 18410 30760 18450 30790
rect 17470 30720 18450 30760
rect 17470 30640 17510 30720
rect 17250 30600 17510 30640
rect 17860 30610 18860 30650
rect 17860 30310 17920 30610
rect 18220 30480 18330 30610
rect 18220 30400 18240 30480
rect 18310 30400 18330 30480
rect 18220 30390 18330 30400
rect 18800 30310 18860 30610
rect 19850 30600 19900 30830
rect 19990 30750 20090 30770
rect 19990 30690 20010 30750
rect 20070 30690 20090 30750
rect 20130 30760 20190 30770
rect 20130 30750 20340 30760
rect 20130 30710 20140 30750
rect 20180 30710 20280 30750
rect 20320 30710 20340 30750
rect 20130 30700 20340 30710
rect 20130 30690 20190 30700
rect 19990 30670 20090 30690
rect 20010 30600 20090 30610
rect 19850 30560 20030 30600
rect 20070 30560 20090 30600
rect 20010 30550 20090 30560
rect 20560 30480 20620 31180
rect 20960 30900 21060 30920
rect 20720 30840 20820 30860
rect 20720 30760 20740 30840
rect 20800 30760 20820 30840
rect 20960 30840 20980 30900
rect 21040 30840 21060 30900
rect 20960 30820 21060 30840
rect 21200 30890 21300 30910
rect 21390 30890 21430 31380
rect 21470 31370 21550 31380
rect 22140 31420 22220 31430
rect 22580 31420 22800 31430
rect 22140 31380 22160 31420
rect 22200 31380 22310 31420
rect 22140 31370 22220 31380
rect 22270 31320 22310 31380
rect 22580 31380 22600 31420
rect 22640 31380 22740 31420
rect 22780 31380 22800 31420
rect 22580 31370 22800 31380
rect 23040 31420 23120 31430
rect 23040 31380 23060 31420
rect 23100 31380 23120 31420
rect 23040 31370 23120 31380
rect 23520 31420 23740 31430
rect 23520 31380 23540 31420
rect 23580 31380 23680 31420
rect 23720 31380 23740 31420
rect 23520 31370 23740 31380
rect 23980 31420 24060 31430
rect 24970 31420 25050 31430
rect 23980 31380 24000 31420
rect 24040 31380 24060 31420
rect 23980 31370 24060 31380
rect 24810 31380 24990 31420
rect 25030 31380 25050 31420
rect 25090 31410 25240 31450
rect 25280 31410 25300 31450
rect 25090 31400 25300 31410
rect 22240 31300 22350 31320
rect 22240 31230 22260 31300
rect 22330 31230 22350 31300
rect 22660 31290 22720 31370
rect 22660 31250 22670 31290
rect 22710 31250 22720 31290
rect 22660 31230 22720 31250
rect 23600 31290 23660 31370
rect 23600 31250 23610 31290
rect 23650 31250 23660 31290
rect 23600 31230 23660 31250
rect 22240 31210 22350 31230
rect 21200 30850 21250 30890
rect 21290 30850 21430 30890
rect 21200 30830 21300 30850
rect 20720 30740 20820 30760
rect 20740 30480 20800 30740
rect 22270 30630 22310 31210
rect 23240 31170 23640 31200
rect 23240 31160 23650 31170
rect 22870 31130 22950 31140
rect 23240 31130 23290 31160
rect 22870 31090 22890 31130
rect 22930 31090 23290 31130
rect 23560 31150 23650 31160
rect 22870 31080 22950 31090
rect 23560 31080 23570 31150
rect 23640 31080 23650 31150
rect 23560 31060 23650 31080
rect 22470 30830 22550 30840
rect 22470 30790 22490 30830
rect 22530 30790 22550 30830
rect 22470 30780 22550 30790
rect 23410 30830 23490 30840
rect 23410 30790 23430 30830
rect 23470 30790 23490 30830
rect 23590 30830 23640 31060
rect 24810 30900 24860 31380
rect 24970 31370 25050 31380
rect 25340 31300 26060 31320
rect 25340 31260 25430 31300
rect 25470 31260 26060 31300
rect 25340 31240 26060 31260
rect 23990 30880 24220 30900
rect 24330 30880 24390 30900
rect 23990 30840 24150 30880
rect 24190 30840 24340 30880
rect 24380 30840 24390 30880
rect 23700 30830 23780 30840
rect 23590 30790 23720 30830
rect 23760 30790 23780 30830
rect 23990 30820 24220 30840
rect 24330 30820 24390 30840
rect 24430 30880 24540 30900
rect 24590 30880 24650 30900
rect 24430 30840 24490 30880
rect 24530 30840 24600 30880
rect 24640 30840 24650 30880
rect 24430 30820 24540 30840
rect 24590 30820 24650 30840
rect 24690 30880 24860 30900
rect 24690 30840 24740 30880
rect 24780 30840 24860 30880
rect 24690 30820 24860 30840
rect 23410 30780 23490 30790
rect 23700 30780 23780 30790
rect 22490 30750 22530 30780
rect 23430 30750 23470 30780
rect 22490 30710 23470 30750
rect 22490 30630 22530 30710
rect 22270 30590 22530 30630
rect 22880 30610 23880 30650
rect 20540 30460 20640 30480
rect 20540 30380 20560 30460
rect 20620 30380 20640 30460
rect 20540 30360 20640 30380
rect 20720 30460 20820 30480
rect 20720 30380 20740 30460
rect 20800 30380 20820 30460
rect 20720 30360 20820 30380
rect 17670 30300 18100 30310
rect 17670 30260 17690 30300
rect 17730 30260 17870 30300
rect 17910 30260 18040 30300
rect 18080 30260 18100 30300
rect 17670 30250 18100 30260
rect 18610 30300 19040 30310
rect 22880 30300 22940 30610
rect 23240 30480 23340 30610
rect 23240 30400 23260 30480
rect 23320 30400 23340 30480
rect 23240 30390 23340 30400
rect 23820 30300 23880 30610
rect 24810 30590 24860 30820
rect 24950 30740 25050 30760
rect 24950 30680 24970 30740
rect 25030 30680 25050 30740
rect 25090 30750 25150 30760
rect 25090 30740 25300 30750
rect 25090 30700 25100 30740
rect 25140 30700 25240 30740
rect 25280 30700 25300 30740
rect 25090 30690 25300 30700
rect 25090 30680 25150 30690
rect 24950 30660 25050 30680
rect 24970 30590 25050 30600
rect 24810 30550 24990 30590
rect 25030 30550 25050 30590
rect 24970 30540 25050 30550
rect 18610 30260 18630 30300
rect 18670 30260 18810 30300
rect 18850 30260 18980 30300
rect 19020 30260 19040 30300
rect 18610 30250 19040 30260
rect 22690 30290 23120 30300
rect 22690 30250 22710 30290
rect 22750 30250 22890 30290
rect 22930 30250 23060 30290
rect 23100 30250 23120 30290
rect 22690 30240 23120 30250
rect 23630 30290 24060 30300
rect 23630 30250 23650 30290
rect 23690 30250 23830 30290
rect 23870 30250 24000 30290
rect 24040 30250 24060 30290
rect 23630 30240 24060 30250
rect 14830 30130 25680 30140
rect 14830 30060 14870 30130
rect 14930 30060 14970 30130
rect 15030 30060 15070 30130
rect 15130 30060 15170 30130
rect 15230 30060 15270 30130
rect 15330 30060 15370 30130
rect 15430 30060 15470 30130
rect 15530 30060 15570 30130
rect 15630 30060 15670 30130
rect 15730 30060 15780 30130
rect 15840 30060 15880 30130
rect 15940 30060 15990 30130
rect 16050 30060 16130 30130
rect 16190 30060 16270 30130
rect 16330 30060 16370 30130
rect 16430 30060 16470 30130
rect 16530 30060 16570 30130
rect 16630 30060 16670 30130
rect 16730 30060 16770 30130
rect 16830 30060 16870 30130
rect 16930 30060 16970 30130
rect 17030 30060 17070 30130
rect 17130 30060 17170 30130
rect 17230 30060 17270 30130
rect 17330 30060 17370 30130
rect 17430 30060 17470 30130
rect 17530 30060 17570 30130
rect 17630 30060 17670 30130
rect 17730 30060 17770 30130
rect 17830 30060 17870 30130
rect 17930 30060 17970 30130
rect 18030 30060 18070 30130
rect 18130 30060 18170 30130
rect 18230 30060 18270 30130
rect 18330 30060 18370 30130
rect 18430 30060 18470 30130
rect 18530 30060 18570 30130
rect 18630 30060 18670 30130
rect 18730 30060 18770 30130
rect 18830 30060 18870 30130
rect 18930 30060 18970 30130
rect 19030 30060 19070 30130
rect 19130 30060 19170 30130
rect 19230 30060 19270 30130
rect 19330 30060 19370 30130
rect 19430 30060 19470 30130
rect 19530 30060 19570 30130
rect 19630 30060 19670 30130
rect 19730 30060 19770 30130
rect 19830 30060 19870 30130
rect 19930 30060 19970 30130
rect 20030 30060 20070 30130
rect 20130 30060 20170 30130
rect 20230 30060 20270 30130
rect 20330 30060 20370 30130
rect 20430 30060 20470 30130
rect 20530 30060 20570 30130
rect 20630 30060 20670 30130
rect 20730 30060 20770 30130
rect 20830 30060 20870 30130
rect 20930 30060 20970 30130
rect 21030 30060 21070 30130
rect 21130 30060 21170 30130
rect 21230 30060 21270 30130
rect 21330 30060 21370 30130
rect 21430 30060 21470 30130
rect 21530 30060 21570 30130
rect 21630 30060 21670 30130
rect 21730 30060 21770 30130
rect 21830 30060 21870 30130
rect 21930 30060 21970 30130
rect 22030 30060 22070 30130
rect 22130 30060 22170 30130
rect 22230 30060 22270 30130
rect 22330 30060 22370 30130
rect 22430 30060 22470 30130
rect 22530 30060 22570 30130
rect 22630 30060 22670 30130
rect 22730 30060 22770 30130
rect 22830 30060 22870 30130
rect 22930 30060 22970 30130
rect 23030 30060 23070 30130
rect 23130 30060 23170 30130
rect 23230 30060 23270 30130
rect 23330 30060 23370 30130
rect 23430 30060 23470 30130
rect 23530 30060 23570 30130
rect 23630 30060 23670 30130
rect 23730 30060 23770 30130
rect 23830 30060 23870 30130
rect 23930 30060 23970 30130
rect 24030 30060 24070 30130
rect 24130 30060 24170 30130
rect 24230 30060 24270 30130
rect 24330 30060 24370 30130
rect 24430 30060 24470 30130
rect 24530 30060 24570 30130
rect 24630 30060 24670 30130
rect 24730 30060 24770 30130
rect 24830 30060 24870 30130
rect 24930 30060 24970 30130
rect 25030 30060 25070 30130
rect 25130 30060 25170 30130
rect 25230 30060 25270 30130
rect 25330 30060 25370 30130
rect 25430 30060 25470 30130
rect 25530 30060 25570 30130
rect 25630 30060 25680 30130
rect 14830 29980 25680 30060
rect 14830 29170 22440 29980
rect 23080 29170 25680 29980
rect 14830 29120 25680 29170
rect 22390 29110 23130 29120
rect 12700 28620 12840 28640
rect 25970 28620 26060 31240
rect 12700 28510 12720 28620
rect 12820 28510 26060 28620
rect 12700 28490 12840 28510
rect 12690 28270 12830 28290
rect 26320 28270 26430 35310
rect 12690 28160 12710 28270
rect 12810 28160 26430 28270
rect 12690 28140 12830 28160
rect 6910 27810 11690 27910
rect 6910 25480 7000 27810
rect 7320 27360 20640 27430
rect 7320 26670 7370 27360
rect 8200 26670 8400 27360
rect 9230 26670 9430 27360
rect 10260 26670 10460 27360
rect 11290 26670 11490 27360
rect 12320 26670 12520 27360
rect 13350 26670 13550 27360
rect 14380 26670 14580 27360
rect 15410 26670 15610 27360
rect 16440 26670 16640 27360
rect 17470 26670 17670 27360
rect 18500 26670 18700 27360
rect 19530 26670 19760 27360
rect 20590 26670 20640 27360
rect 7320 26610 20640 26670
rect 7320 26570 7360 26610
rect 7400 26570 7440 26610
rect 7480 26570 7520 26610
rect 7560 26570 7600 26610
rect 7640 26570 7680 26610
rect 7720 26570 7760 26610
rect 7800 26570 7840 26610
rect 7880 26570 7920 26610
rect 7960 26570 8000 26610
rect 8040 26570 8080 26610
rect 8120 26570 8160 26610
rect 8200 26570 8240 26610
rect 8280 26570 8320 26610
rect 8360 26570 8400 26610
rect 8440 26570 8480 26610
rect 8520 26570 8560 26610
rect 8600 26570 8640 26610
rect 8680 26570 8720 26610
rect 8760 26570 8800 26610
rect 8840 26570 8880 26610
rect 8920 26570 8960 26610
rect 9000 26570 9040 26610
rect 9080 26570 9120 26610
rect 9160 26570 9200 26610
rect 9240 26570 9280 26610
rect 9320 26570 9360 26610
rect 9400 26570 9440 26610
rect 9480 26570 9520 26610
rect 9560 26570 9600 26610
rect 9640 26570 9680 26610
rect 9720 26570 9760 26610
rect 9800 26570 9840 26610
rect 9880 26570 9920 26610
rect 9960 26570 10000 26610
rect 10040 26570 10080 26610
rect 10120 26570 10160 26610
rect 10200 26570 10240 26610
rect 10280 26570 10320 26610
rect 10360 26570 10400 26610
rect 10440 26570 10480 26610
rect 10520 26570 10560 26610
rect 10600 26570 10640 26610
rect 10680 26570 10720 26610
rect 10760 26570 10800 26610
rect 10840 26570 10880 26610
rect 10920 26570 10960 26610
rect 11000 26570 11040 26610
rect 11080 26570 11120 26610
rect 11160 26570 11200 26610
rect 11240 26570 11280 26610
rect 11320 26570 11360 26610
rect 11400 26570 11440 26610
rect 11480 26570 11520 26610
rect 11560 26570 11600 26610
rect 11640 26570 11680 26610
rect 11720 26570 11760 26610
rect 11800 26570 11840 26610
rect 11880 26570 11920 26610
rect 11960 26570 12000 26610
rect 12040 26570 12080 26610
rect 12120 26570 12160 26610
rect 12200 26570 12240 26610
rect 12280 26570 12320 26610
rect 12360 26570 12400 26610
rect 12440 26570 12480 26610
rect 12520 26570 12560 26610
rect 12600 26570 12640 26610
rect 12680 26570 12720 26610
rect 12760 26570 12800 26610
rect 12840 26570 12880 26610
rect 12920 26570 12960 26610
rect 13000 26570 13040 26610
rect 13080 26570 13120 26610
rect 13160 26570 13200 26610
rect 13240 26570 13280 26610
rect 13320 26570 13360 26610
rect 13400 26570 13440 26610
rect 13480 26570 13520 26610
rect 13560 26570 13600 26610
rect 13640 26570 13680 26610
rect 13720 26570 13760 26610
rect 13800 26570 13840 26610
rect 13880 26570 13920 26610
rect 13960 26570 14000 26610
rect 14040 26570 14080 26610
rect 14120 26570 14160 26610
rect 14200 26570 14240 26610
rect 14280 26570 14320 26610
rect 14360 26570 14400 26610
rect 14440 26570 14480 26610
rect 14520 26570 14560 26610
rect 14600 26570 14640 26610
rect 14680 26570 14720 26610
rect 14760 26570 14800 26610
rect 14840 26570 14880 26610
rect 14920 26570 14960 26610
rect 15000 26570 15040 26610
rect 15080 26570 15120 26610
rect 15160 26570 15200 26610
rect 15240 26570 15280 26610
rect 15320 26570 15360 26610
rect 15400 26570 15440 26610
rect 15480 26570 15520 26610
rect 15560 26570 15600 26610
rect 15640 26570 15680 26610
rect 15720 26570 15760 26610
rect 15800 26570 15840 26610
rect 15880 26570 15920 26610
rect 15960 26570 16000 26610
rect 16040 26570 16080 26610
rect 16120 26570 16160 26610
rect 16200 26570 16240 26610
rect 16280 26570 16320 26610
rect 16360 26570 16400 26610
rect 16440 26570 16480 26610
rect 16520 26570 16560 26610
rect 16600 26570 16640 26610
rect 16680 26570 16720 26610
rect 16760 26570 16800 26610
rect 16840 26570 16880 26610
rect 16920 26570 16960 26610
rect 17000 26570 17040 26610
rect 17080 26570 17120 26610
rect 17160 26570 17200 26610
rect 17240 26570 17280 26610
rect 17320 26570 17360 26610
rect 17400 26570 17440 26610
rect 17480 26570 17520 26610
rect 17560 26570 17600 26610
rect 17640 26570 17680 26610
rect 17720 26570 17760 26610
rect 17800 26570 17840 26610
rect 17880 26570 17920 26610
rect 17960 26570 18000 26610
rect 18040 26570 18080 26610
rect 18120 26570 18160 26610
rect 18200 26570 18240 26610
rect 18280 26570 18320 26610
rect 18360 26570 18400 26610
rect 18440 26570 18480 26610
rect 18520 26570 18560 26610
rect 18600 26570 18640 26610
rect 18680 26570 18720 26610
rect 18760 26570 18800 26610
rect 18840 26570 18880 26610
rect 18920 26570 18960 26610
rect 19000 26570 19040 26610
rect 19080 26570 19120 26610
rect 19160 26570 19200 26610
rect 19240 26570 19280 26610
rect 19320 26570 19360 26610
rect 19400 26570 19440 26610
rect 19480 26570 19520 26610
rect 19560 26570 19600 26610
rect 19640 26570 19680 26610
rect 19720 26570 19760 26610
rect 19800 26570 19840 26610
rect 19880 26570 19920 26610
rect 19960 26570 20000 26610
rect 20040 26570 20080 26610
rect 20120 26570 20160 26610
rect 20200 26570 20240 26610
rect 20280 26570 20320 26610
rect 20360 26570 20400 26610
rect 20440 26570 20480 26610
rect 20520 26570 20560 26610
rect 20600 26570 20640 26610
rect 7320 26560 20640 26570
rect 7060 25560 7920 25580
rect 7060 25500 7080 25560
rect 7140 25500 7820 25560
rect 7880 25500 7920 25560
rect 7060 25480 7920 25500
rect 6740 25190 7390 25210
rect 6740 25130 7290 25190
rect 7350 25130 7390 25190
rect 6740 25110 7390 25130
rect 6740 15120 6820 25110
rect 8370 24960 8420 26560
rect 9510 24960 9550 26560
rect 9660 25950 9740 25960
rect 9660 25910 9680 25950
rect 9720 25910 9740 25950
rect 9660 25900 9740 25910
rect 9920 25950 10000 25960
rect 9920 25910 9940 25950
rect 9980 25910 10000 25950
rect 9920 25900 10000 25910
rect 10650 25950 10730 25960
rect 10650 25910 10670 25950
rect 10710 25910 10730 25950
rect 10650 25900 10730 25910
rect 10910 25950 10990 25960
rect 10910 25910 10930 25950
rect 10970 25910 10990 25950
rect 10910 25900 10990 25910
rect 11650 25950 11730 25960
rect 11650 25910 11670 25950
rect 11710 25910 11730 25950
rect 11650 25900 11730 25910
rect 11910 25950 11990 25960
rect 11910 25910 11930 25950
rect 11970 25910 11990 25950
rect 14110 25950 14190 25960
rect 11910 25900 11990 25910
rect 13210 25930 13290 25940
rect 9680 25070 9720 25900
rect 9940 25070 9980 25900
rect 10670 25070 10710 25900
rect 10930 25070 10970 25900
rect 11670 25070 11710 25900
rect 11930 25070 11970 25900
rect 13210 25890 13230 25930
rect 13270 25890 13290 25930
rect 13210 25880 13290 25890
rect 13550 25930 13630 25940
rect 13550 25890 13570 25930
rect 13610 25890 13630 25930
rect 13550 25880 13630 25890
rect 13770 25930 13850 25940
rect 13770 25890 13790 25930
rect 13830 25890 13850 25930
rect 14110 25910 14130 25950
rect 14170 25910 14190 25950
rect 14110 25900 14190 25910
rect 14330 25950 14410 25960
rect 14330 25910 14350 25950
rect 14390 25910 14410 25950
rect 14330 25900 14410 25910
rect 14550 25950 14630 25960
rect 14550 25910 14570 25950
rect 14610 25910 14630 25950
rect 14550 25900 14630 25910
rect 14770 25950 14850 25960
rect 14770 25910 14790 25950
rect 14830 25910 14850 25950
rect 14770 25900 14850 25910
rect 15170 25950 15250 25960
rect 15170 25910 15190 25950
rect 15230 25910 15250 25950
rect 15170 25900 15250 25910
rect 15390 25950 15470 25960
rect 15390 25910 15410 25950
rect 15450 25910 15470 25950
rect 15390 25900 15470 25910
rect 15610 25950 15690 25960
rect 15610 25910 15630 25950
rect 15670 25910 15690 25950
rect 15610 25900 15690 25910
rect 15830 25950 15910 25960
rect 15830 25910 15850 25950
rect 15890 25910 15910 25950
rect 15830 25900 15910 25910
rect 16050 25950 16130 25960
rect 16050 25910 16070 25950
rect 16110 25910 16130 25950
rect 16050 25900 16130 25910
rect 16270 25950 16350 25960
rect 16270 25910 16290 25950
rect 16330 25910 16350 25950
rect 16270 25900 16350 25910
rect 16490 25950 16570 25960
rect 16490 25910 16510 25950
rect 16550 25910 16570 25950
rect 16490 25900 16570 25910
rect 16710 25950 16790 25960
rect 16710 25910 16730 25950
rect 16770 25910 16790 25950
rect 16710 25900 16790 25910
rect 17120 25950 17200 25960
rect 17120 25910 17140 25950
rect 17180 25910 17200 25950
rect 17120 25900 17200 25910
rect 17340 25950 17420 25960
rect 17340 25910 17360 25950
rect 17400 25910 17420 25950
rect 17340 25900 17420 25910
rect 17560 25950 17640 25960
rect 17560 25910 17580 25950
rect 17620 25910 17640 25950
rect 17560 25900 17640 25910
rect 17780 25950 17860 25960
rect 17780 25910 17800 25950
rect 17840 25910 17860 25950
rect 17780 25900 17860 25910
rect 18000 25950 18080 25960
rect 18000 25910 18020 25950
rect 18060 25910 18080 25950
rect 18000 25900 18080 25910
rect 18220 25950 18300 25960
rect 18220 25910 18240 25950
rect 18280 25910 18300 25950
rect 18220 25900 18300 25910
rect 18440 25950 18520 25960
rect 18440 25910 18460 25950
rect 18500 25910 18520 25950
rect 18440 25900 18520 25910
rect 18660 25950 18740 25960
rect 18660 25910 18680 25950
rect 18720 25910 18740 25950
rect 18660 25900 18740 25910
rect 18880 25950 18960 25960
rect 18880 25910 18900 25950
rect 18940 25910 18960 25950
rect 18880 25900 18960 25910
rect 19100 25950 19180 25960
rect 19100 25910 19120 25950
rect 19160 25910 19180 25950
rect 19100 25900 19180 25910
rect 19320 25950 19400 25960
rect 19320 25910 19340 25950
rect 19380 25910 19400 25950
rect 19320 25900 19400 25910
rect 19540 25950 19620 25960
rect 19540 25910 19560 25950
rect 19600 25910 19620 25950
rect 19540 25900 19620 25910
rect 19760 25950 19840 25960
rect 19760 25910 19780 25950
rect 19820 25910 19840 25950
rect 19760 25900 19840 25910
rect 19980 25950 20060 25960
rect 19980 25910 20000 25950
rect 20040 25910 20060 25950
rect 19980 25900 20060 25910
rect 20200 25950 20280 25960
rect 20200 25910 20220 25950
rect 20260 25910 20280 25950
rect 20200 25900 20280 25910
rect 20420 25950 20500 25960
rect 20420 25910 20440 25950
rect 20480 25910 20500 25950
rect 20420 25900 20500 25910
rect 13770 25880 13850 25890
rect 9660 25060 9740 25070
rect 9660 25020 9680 25060
rect 9720 25020 9740 25060
rect 9660 25010 9740 25020
rect 9920 25060 10000 25070
rect 9920 25020 9940 25060
rect 9980 25020 10000 25060
rect 9920 25010 10000 25020
rect 10650 25060 10730 25070
rect 10650 25020 10670 25060
rect 10710 25020 10730 25060
rect 10650 25010 10730 25020
rect 10910 25060 10990 25070
rect 10910 25020 10930 25060
rect 10970 25020 10990 25060
rect 10910 25010 10990 25020
rect 11650 25060 11730 25070
rect 11650 25020 11670 25060
rect 11710 25020 11730 25060
rect 11650 25010 11730 25020
rect 11910 25060 11990 25070
rect 11910 25020 11930 25060
rect 11970 25020 11990 25060
rect 13230 25050 13270 25880
rect 13570 25050 13610 25880
rect 13790 25050 13830 25880
rect 14130 25070 14170 25900
rect 14350 25070 14390 25900
rect 14570 25070 14610 25900
rect 14790 25070 14830 25900
rect 15190 25070 15230 25900
rect 15410 25070 15450 25900
rect 15630 25070 15670 25900
rect 15850 25070 15890 25900
rect 16070 25070 16110 25900
rect 16290 25070 16330 25900
rect 16510 25070 16550 25900
rect 16730 25070 16770 25900
rect 17140 25070 17180 25900
rect 17360 25070 17400 25900
rect 17580 25070 17620 25900
rect 17800 25070 17840 25900
rect 18020 25070 18060 25900
rect 18240 25070 18280 25900
rect 18460 25070 18500 25900
rect 18680 25070 18720 25900
rect 18900 25070 18940 25900
rect 19120 25070 19160 25900
rect 19340 25070 19380 25900
rect 19560 25070 19600 25900
rect 19780 25070 19820 25900
rect 20000 25070 20040 25900
rect 20220 25070 20260 25900
rect 20440 25070 20480 25900
rect 14110 25060 14190 25070
rect 11910 25010 11990 25020
rect 13210 25040 13290 25050
rect 13210 25000 13230 25040
rect 13270 25000 13290 25040
rect 13210 24990 13290 25000
rect 13550 25040 13630 25050
rect 13550 25000 13570 25040
rect 13610 25000 13630 25040
rect 13550 24990 13630 25000
rect 13770 25040 13850 25050
rect 13770 25000 13790 25040
rect 13830 25000 13850 25040
rect 14110 25020 14130 25060
rect 14170 25020 14190 25060
rect 14110 25010 14190 25020
rect 14330 25060 14410 25070
rect 14330 25020 14350 25060
rect 14390 25020 14410 25060
rect 14330 25010 14410 25020
rect 14550 25060 14630 25070
rect 14550 25020 14570 25060
rect 14610 25020 14630 25060
rect 14550 25010 14630 25020
rect 14770 25060 14850 25070
rect 14770 25020 14790 25060
rect 14830 25020 14850 25060
rect 14770 25010 14850 25020
rect 15170 25060 15250 25070
rect 15170 25020 15190 25060
rect 15230 25020 15250 25060
rect 15170 25010 15250 25020
rect 15390 25060 15470 25070
rect 15390 25020 15410 25060
rect 15450 25020 15470 25060
rect 15390 25010 15470 25020
rect 15610 25060 15690 25070
rect 15610 25020 15630 25060
rect 15670 25020 15690 25060
rect 15610 25010 15690 25020
rect 15830 25060 15910 25070
rect 15830 25020 15850 25060
rect 15890 25020 15910 25060
rect 15830 25010 15910 25020
rect 16050 25060 16130 25070
rect 16050 25020 16070 25060
rect 16110 25020 16130 25060
rect 16050 25010 16130 25020
rect 16270 25060 16350 25070
rect 16270 25020 16290 25060
rect 16330 25020 16350 25060
rect 16270 25010 16350 25020
rect 16490 25060 16570 25070
rect 16490 25020 16510 25060
rect 16550 25020 16570 25060
rect 16490 25010 16570 25020
rect 16710 25060 16790 25070
rect 16710 25020 16730 25060
rect 16770 25020 16790 25060
rect 16710 25010 16790 25020
rect 17120 25060 17200 25070
rect 17120 25020 17140 25060
rect 17180 25020 17200 25060
rect 17120 25010 17200 25020
rect 17340 25060 17420 25070
rect 17340 25020 17360 25060
rect 17400 25020 17420 25060
rect 17340 25010 17420 25020
rect 17560 25060 17640 25070
rect 17560 25020 17580 25060
rect 17620 25020 17640 25060
rect 17560 25010 17640 25020
rect 17780 25060 17860 25070
rect 17780 25020 17800 25060
rect 17840 25020 17860 25060
rect 17780 25010 17860 25020
rect 18000 25060 18080 25070
rect 18000 25020 18020 25060
rect 18060 25020 18080 25060
rect 18000 25010 18080 25020
rect 18220 25060 18300 25070
rect 18220 25020 18240 25060
rect 18280 25020 18300 25060
rect 18220 25010 18300 25020
rect 18440 25060 18520 25070
rect 18440 25020 18460 25060
rect 18500 25020 18520 25060
rect 18440 25010 18520 25020
rect 18660 25060 18740 25070
rect 18660 25020 18680 25060
rect 18720 25020 18740 25060
rect 18660 25010 18740 25020
rect 18880 25060 18960 25070
rect 18880 25020 18900 25060
rect 18940 25020 18960 25060
rect 18880 25010 18960 25020
rect 19100 25060 19180 25070
rect 19100 25020 19120 25060
rect 19160 25020 19180 25060
rect 19100 25010 19180 25020
rect 19320 25060 19400 25070
rect 19320 25020 19340 25060
rect 19380 25020 19400 25060
rect 19320 25010 19400 25020
rect 19540 25060 19620 25070
rect 19540 25020 19560 25060
rect 19600 25020 19620 25060
rect 19540 25010 19620 25020
rect 19760 25060 19840 25070
rect 19760 25020 19780 25060
rect 19820 25020 19840 25060
rect 19760 25010 19840 25020
rect 19980 25060 20060 25070
rect 19980 25020 20000 25060
rect 20040 25020 20060 25060
rect 19980 25010 20060 25020
rect 20200 25060 20280 25070
rect 20200 25020 20220 25060
rect 20260 25020 20280 25060
rect 20200 25010 20280 25020
rect 20420 25060 20500 25070
rect 20420 25020 20440 25060
rect 20480 25020 20500 25060
rect 20420 25010 20500 25020
rect 13770 24990 13850 25000
rect 8370 24940 8550 24960
rect 8370 24900 8500 24940
rect 8540 24900 8550 24940
rect 8730 24940 8930 24960
rect 8730 24920 8800 24940
rect 8480 24880 8550 24900
rect 8740 24900 8800 24920
rect 8840 24900 8880 24940
rect 8920 24900 8930 24940
rect 8740 24880 8930 24900
rect 8970 24950 9070 24960
rect 8970 24890 8990 24950
rect 9050 24890 9070 24950
rect 9200 24950 9290 24960
rect 9200 24910 9220 24950
rect 9260 24910 9290 24950
rect 9200 24900 9290 24910
rect 9510 24940 9630 24960
rect 9510 24900 9580 24940
rect 9620 24900 9630 24940
rect 9930 24950 10230 24960
rect 9930 24910 10080 24950
rect 10120 24910 10160 24950
rect 10200 24910 10230 24950
rect 9930 24900 10230 24910
rect 10340 24950 10620 24960
rect 10340 24910 10460 24950
rect 10500 24940 10620 24950
rect 10500 24910 10570 24940
rect 10340 24900 10570 24910
rect 10610 24900 10620 24940
rect 10920 24950 11220 24960
rect 10920 24910 11070 24950
rect 11110 24910 11150 24950
rect 11190 24910 11220 24950
rect 10920 24900 11220 24910
rect 11330 24950 11620 24960
rect 11330 24910 11450 24950
rect 11490 24940 11620 24950
rect 11490 24910 11570 24940
rect 11330 24900 11570 24910
rect 11610 24900 11620 24940
rect 11920 24950 12220 24960
rect 11920 24910 12070 24950
rect 12110 24910 12150 24950
rect 12190 24910 12220 24950
rect 11920 24900 12220 24910
rect 12330 24950 12600 24960
rect 12330 24910 12450 24950
rect 12490 24910 12530 24950
rect 12570 24910 12600 24950
rect 12330 24900 12600 24910
rect 12710 24940 12950 24960
rect 12710 24900 12820 24940
rect 12860 24900 12900 24940
rect 12940 24900 12950 24940
rect 8970 24880 9070 24890
rect 8060 24870 8160 24880
rect 8060 24860 8080 24870
rect 8030 24800 8080 24860
rect 8140 24850 8160 24870
rect 8630 24860 8700 24880
rect 8740 24870 8800 24880
rect 8630 24850 8650 24860
rect 8140 24820 8650 24850
rect 8690 24820 8700 24860
rect 8140 24800 8700 24820
rect 8060 24790 8160 24800
rect 7530 24770 7650 24790
rect 7500 24710 7570 24770
rect 7630 24710 7650 24770
rect 8180 24730 8280 24750
rect 9210 24730 9260 24900
rect 9510 24880 9630 24900
rect 10560 24880 10620 24900
rect 11560 24880 11620 24900
rect 12710 24880 12950 24900
rect 12990 24940 13180 24960
rect 12990 24900 13000 24940
rect 13040 24900 13130 24940
rect 13170 24900 13180 24940
rect 12990 24880 13180 24900
rect 13330 24940 13520 24960
rect 13330 24900 13340 24940
rect 13380 24900 13470 24940
rect 13510 24900 13520 24940
rect 13330 24880 13520 24900
rect 13890 24940 14080 24960
rect 13890 24900 13900 24940
rect 13940 24900 14030 24940
rect 14070 24900 14080 24940
rect 13890 24880 14080 24900
rect 14890 24940 15140 24960
rect 14890 24900 14900 24940
rect 14940 24900 15090 24940
rect 15130 24900 15140 24940
rect 14890 24880 15140 24900
rect 16830 24940 16960 24950
rect 17020 24940 17090 24960
rect 16830 24890 16890 24940
rect 16940 24900 17040 24940
rect 17080 24900 17090 24940
rect 16940 24890 16960 24900
rect 16830 24880 16960 24890
rect 17020 24880 17090 24900
rect 20540 24940 23510 24950
rect 20540 24890 20600 24940
rect 20650 24890 23510 24940
rect 20540 24880 23510 24890
rect 9830 24840 9890 24860
rect 9400 24800 9840 24840
rect 9880 24800 9890 24840
rect 9830 24780 9890 24800
rect 10400 24850 10490 24870
rect 10400 24790 10410 24850
rect 10480 24840 10490 24850
rect 10820 24840 10880 24860
rect 10480 24800 10830 24840
rect 10870 24800 10880 24840
rect 10480 24790 10490 24800
rect 10400 24770 10490 24790
rect 10820 24780 10880 24800
rect 11400 24850 11490 24870
rect 11400 24790 11410 24850
rect 11480 24840 11490 24850
rect 11820 24840 11880 24860
rect 11480 24800 11830 24840
rect 11870 24800 11880 24840
rect 11480 24790 11490 24800
rect 11400 24770 11490 24790
rect 11820 24780 11880 24800
rect 7530 24690 7650 24710
rect 8170 24670 8200 24730
rect 8260 24670 9260 24730
rect 8180 24650 8280 24670
rect 9080 24610 9170 24630
rect 9080 24560 9100 24610
rect 9150 24560 9170 24610
rect 9080 24540 9170 24560
rect 9090 24460 9160 24540
rect 9080 24440 9170 24460
rect 9080 24380 9090 24440
rect 9160 24380 9170 24440
rect 9080 24360 9170 24380
rect 7280 24290 20620 24300
rect 7280 24250 7320 24290
rect 7360 24250 7400 24290
rect 7440 24250 7480 24290
rect 7520 24250 7560 24290
rect 7600 24250 7640 24290
rect 7680 24250 7720 24290
rect 7760 24250 7800 24290
rect 7840 24250 7890 24290
rect 7930 24250 7970 24290
rect 8010 24250 8050 24290
rect 8090 24250 8130 24290
rect 8170 24250 8210 24290
rect 8250 24250 8290 24290
rect 8330 24250 8400 24290
rect 8440 24250 8520 24290
rect 8560 24250 8600 24290
rect 8640 24250 8680 24290
rect 8720 24250 8760 24290
rect 8800 24250 8840 24290
rect 8880 24250 8920 24290
rect 8960 24250 9000 24290
rect 9040 24250 9080 24290
rect 9120 24250 9160 24290
rect 9200 24250 9270 24290
rect 9310 24250 9350 24290
rect 9390 24250 9430 24290
rect 9470 24250 9510 24290
rect 9550 24250 9590 24290
rect 9630 24250 9670 24290
rect 9710 24250 9750 24290
rect 9790 24250 9830 24290
rect 9870 24250 9910 24290
rect 9950 24250 9990 24290
rect 10030 24250 10070 24290
rect 10110 24250 10150 24290
rect 10190 24250 10230 24290
rect 10270 24250 10310 24290
rect 10350 24250 10390 24290
rect 10430 24250 10470 24290
rect 10510 24250 10550 24290
rect 10590 24250 10630 24290
rect 10670 24250 10710 24290
rect 10750 24250 10790 24290
rect 10830 24250 10870 24290
rect 10910 24250 10950 24290
rect 10990 24250 11030 24290
rect 11070 24250 11110 24290
rect 11150 24250 11190 24290
rect 11230 24250 11270 24290
rect 11310 24250 11350 24290
rect 11390 24250 11430 24290
rect 11470 24250 11510 24290
rect 11550 24250 11590 24290
rect 11630 24250 11670 24290
rect 11710 24250 11750 24290
rect 11790 24250 11830 24290
rect 11870 24250 11910 24290
rect 11950 24250 11990 24290
rect 12030 24250 12070 24290
rect 12110 24250 12150 24290
rect 12190 24250 12230 24290
rect 12270 24250 12310 24290
rect 12350 24250 12390 24290
rect 12430 24250 12470 24290
rect 12510 24250 12550 24290
rect 12590 24250 12630 24290
rect 12670 24250 12710 24290
rect 12750 24250 12790 24290
rect 12830 24250 12870 24290
rect 12910 24250 12950 24290
rect 12990 24250 13030 24290
rect 13070 24250 13110 24290
rect 13150 24250 13190 24290
rect 13230 24250 13270 24290
rect 13310 24250 13350 24290
rect 13390 24250 13430 24290
rect 13470 24250 13510 24290
rect 13550 24250 13590 24290
rect 13630 24250 13670 24290
rect 13710 24250 13750 24290
rect 13790 24250 13830 24290
rect 13870 24250 13910 24290
rect 13950 24250 13990 24290
rect 14030 24250 14070 24290
rect 14110 24250 14150 24290
rect 14190 24250 14230 24290
rect 14270 24250 14310 24290
rect 14350 24250 14390 24290
rect 14430 24250 14470 24290
rect 14510 24250 14550 24290
rect 14590 24250 14630 24290
rect 14670 24250 14710 24290
rect 14750 24250 14790 24290
rect 14830 24250 14870 24290
rect 14910 24250 14950 24290
rect 14990 24250 15030 24290
rect 15070 24250 15110 24290
rect 15150 24250 15190 24290
rect 15230 24250 15270 24290
rect 15310 24250 15350 24290
rect 15390 24250 15430 24290
rect 15470 24250 15510 24290
rect 15550 24250 15590 24290
rect 15630 24250 15670 24290
rect 15710 24250 15750 24290
rect 15790 24250 15830 24290
rect 15870 24250 15910 24290
rect 15950 24250 15990 24290
rect 16030 24250 16070 24290
rect 16110 24250 16150 24290
rect 16190 24250 16230 24290
rect 16270 24250 16310 24290
rect 16350 24250 16390 24290
rect 16430 24250 16470 24290
rect 16510 24250 16550 24290
rect 16590 24250 16630 24290
rect 16670 24250 16710 24290
rect 16750 24250 16790 24290
rect 16830 24250 16870 24290
rect 16910 24250 16950 24290
rect 16990 24250 17030 24290
rect 17070 24250 17110 24290
rect 17150 24250 17190 24290
rect 17230 24250 17270 24290
rect 17310 24250 17350 24290
rect 17390 24250 17430 24290
rect 17470 24250 17510 24290
rect 17550 24250 17590 24290
rect 17630 24250 17670 24290
rect 17710 24250 17750 24290
rect 17790 24250 17830 24290
rect 17870 24250 17910 24290
rect 17950 24250 17990 24290
rect 18030 24250 18070 24290
rect 18110 24250 18150 24290
rect 18190 24250 18230 24290
rect 18270 24250 18310 24290
rect 18350 24250 18390 24290
rect 18430 24250 18470 24290
rect 18510 24250 18550 24290
rect 18590 24250 18630 24290
rect 18670 24250 18710 24290
rect 18750 24250 18790 24290
rect 18830 24250 18870 24290
rect 18910 24250 18950 24290
rect 18990 24250 19030 24290
rect 19070 24250 19110 24290
rect 19150 24250 19190 24290
rect 19230 24250 19270 24290
rect 19310 24250 19350 24290
rect 19390 24250 19430 24290
rect 19470 24250 19510 24290
rect 19550 24250 19590 24290
rect 19630 24250 19670 24290
rect 19710 24250 19750 24290
rect 19790 24250 19830 24290
rect 19870 24250 19910 24290
rect 19950 24250 19990 24290
rect 20030 24250 20070 24290
rect 20110 24250 20150 24290
rect 20190 24250 20230 24290
rect 20270 24250 20310 24290
rect 20350 24250 20390 24290
rect 20430 24250 20470 24290
rect 20510 24250 20550 24290
rect 20590 24250 20620 24290
rect 7280 24190 20620 24250
rect 7280 23380 19560 24190
rect 20370 23380 20620 24190
rect 7280 23320 20620 23380
rect 7280 23280 7310 23320
rect 7350 23280 7390 23320
rect 7430 23280 7470 23320
rect 7510 23280 7550 23320
rect 7590 23280 7630 23320
rect 7670 23280 7710 23320
rect 7750 23280 7790 23320
rect 7830 23280 7870 23320
rect 7910 23280 7950 23320
rect 7990 23280 8030 23320
rect 8070 23280 8110 23320
rect 8150 23280 8190 23320
rect 8230 23280 8270 23320
rect 8310 23280 8350 23320
rect 8390 23280 8430 23320
rect 8470 23280 8520 23320
rect 8560 23280 8600 23320
rect 8640 23280 8680 23320
rect 8720 23280 8760 23320
rect 8800 23280 8840 23320
rect 8880 23280 8920 23320
rect 8960 23280 9000 23320
rect 9040 23280 9080 23320
rect 9120 23280 9160 23320
rect 9200 23280 9270 23320
rect 9310 23280 9350 23320
rect 9390 23280 9430 23320
rect 9470 23280 9510 23320
rect 9550 23280 9590 23320
rect 9630 23280 9670 23320
rect 9710 23280 9750 23320
rect 9790 23280 9830 23320
rect 9870 23280 9910 23320
rect 9950 23280 9990 23320
rect 10030 23280 10070 23320
rect 10110 23280 10150 23320
rect 10190 23280 10230 23320
rect 10270 23280 10310 23320
rect 10350 23280 10390 23320
rect 10430 23280 10470 23320
rect 10510 23280 10550 23320
rect 10590 23280 10630 23320
rect 10670 23280 10710 23320
rect 10750 23280 10790 23320
rect 10830 23280 10870 23320
rect 10910 23280 10950 23320
rect 10990 23280 11030 23320
rect 11070 23280 11110 23320
rect 11150 23280 11190 23320
rect 11230 23280 11270 23320
rect 11310 23280 11350 23320
rect 11390 23280 11430 23320
rect 11470 23280 11510 23320
rect 11550 23280 11590 23320
rect 11630 23280 11670 23320
rect 11710 23280 11750 23320
rect 11790 23280 11830 23320
rect 11870 23280 11910 23320
rect 11950 23280 11990 23320
rect 12030 23280 12070 23320
rect 12110 23280 12150 23320
rect 12190 23280 12230 23320
rect 12270 23280 12310 23320
rect 12350 23280 12390 23320
rect 12430 23280 12470 23320
rect 12510 23280 12550 23320
rect 12590 23280 12630 23320
rect 12670 23280 12710 23320
rect 12750 23280 12790 23320
rect 12830 23280 12870 23320
rect 12910 23280 12950 23320
rect 12990 23280 13030 23320
rect 13070 23280 13110 23320
rect 13150 23280 13190 23320
rect 13230 23280 13270 23320
rect 13310 23280 13350 23320
rect 13390 23280 13430 23320
rect 13470 23280 13510 23320
rect 13550 23280 13590 23320
rect 13630 23280 13670 23320
rect 13710 23280 13750 23320
rect 13790 23280 13830 23320
rect 13870 23280 13910 23320
rect 13950 23280 13990 23320
rect 14030 23280 14070 23320
rect 14110 23280 14150 23320
rect 14190 23280 14230 23320
rect 14270 23280 14310 23320
rect 14350 23280 14390 23320
rect 14430 23280 14470 23320
rect 14510 23280 14550 23320
rect 14590 23280 14630 23320
rect 14670 23280 14710 23320
rect 14750 23280 14790 23320
rect 14830 23280 14870 23320
rect 14910 23280 14950 23320
rect 14990 23280 15030 23320
rect 15070 23280 15110 23320
rect 15150 23280 15190 23320
rect 15230 23280 15270 23320
rect 15310 23280 15350 23320
rect 15390 23280 15430 23320
rect 15470 23280 15510 23320
rect 15550 23280 15590 23320
rect 15630 23280 15670 23320
rect 15710 23280 15750 23320
rect 15790 23280 15830 23320
rect 15870 23280 15910 23320
rect 15950 23280 15990 23320
rect 16030 23280 16070 23320
rect 16110 23280 16150 23320
rect 16190 23280 16230 23320
rect 16270 23280 16310 23320
rect 16350 23280 16390 23320
rect 16430 23280 16470 23320
rect 16510 23280 16550 23320
rect 16590 23280 16630 23320
rect 16670 23280 16710 23320
rect 16750 23280 16790 23320
rect 16830 23280 16870 23320
rect 16910 23280 16950 23320
rect 16990 23280 17030 23320
rect 17070 23280 17110 23320
rect 17150 23280 17190 23320
rect 17230 23280 17270 23320
rect 17310 23280 17350 23320
rect 17390 23280 17430 23320
rect 17470 23280 17510 23320
rect 17550 23280 17590 23320
rect 17630 23280 17670 23320
rect 17710 23280 17750 23320
rect 17790 23280 17830 23320
rect 17870 23280 17910 23320
rect 17950 23280 17990 23320
rect 18030 23280 18070 23320
rect 18110 23280 18150 23320
rect 18190 23280 18230 23320
rect 18270 23280 18310 23320
rect 18350 23280 18390 23320
rect 18430 23280 18470 23320
rect 18510 23280 18550 23320
rect 18590 23280 18630 23320
rect 18670 23280 18710 23320
rect 18750 23280 18790 23320
rect 18830 23280 18870 23320
rect 18910 23280 18950 23320
rect 18990 23280 19030 23320
rect 19070 23280 19110 23320
rect 19150 23280 19190 23320
rect 19230 23280 19270 23320
rect 19310 23280 19350 23320
rect 19390 23280 19430 23320
rect 19470 23280 19510 23320
rect 19550 23280 19590 23320
rect 19630 23280 19670 23320
rect 19710 23280 19750 23320
rect 19790 23280 19830 23320
rect 19870 23280 19910 23320
rect 19950 23280 19990 23320
rect 20030 23280 20070 23320
rect 20110 23280 20150 23320
rect 20190 23280 20230 23320
rect 20270 23280 20310 23320
rect 20350 23280 20390 23320
rect 20430 23280 20470 23320
rect 20510 23280 20550 23320
rect 20590 23280 20620 23320
rect 7280 23270 20620 23280
rect 9080 23140 9170 23160
rect 9080 23080 9090 23140
rect 9160 23080 9170 23140
rect 9080 23060 9170 23080
rect 9090 22930 9160 23060
rect 9080 22910 9170 22930
rect 9080 22860 9100 22910
rect 9150 22860 9170 22910
rect 9080 22840 9170 22860
rect 6940 22770 7690 22790
rect 9830 22770 9890 22790
rect 6940 22730 7640 22770
rect 7680 22730 7690 22770
rect 6940 18680 7040 22730
rect 7630 22710 7690 22730
rect 8260 22750 8700 22770
rect 8260 22720 8650 22750
rect 7370 22680 7430 22700
rect 8260 22680 8310 22720
rect 8630 22710 8650 22720
rect 8690 22710 8700 22750
rect 9830 22730 9840 22770
rect 9880 22730 9890 22770
rect 8630 22690 8700 22710
rect 9200 22700 9290 22720
rect 9830 22710 9890 22730
rect 10400 22780 10490 22800
rect 10400 22720 10410 22780
rect 10480 22770 10490 22780
rect 10820 22770 10880 22790
rect 10480 22730 10830 22770
rect 10870 22730 10880 22770
rect 10480 22720 10490 22730
rect 10400 22700 10490 22720
rect 10820 22710 10880 22730
rect 11400 22780 11490 22800
rect 11400 22720 11410 22780
rect 11480 22770 11490 22780
rect 11820 22770 11880 22790
rect 11480 22730 11830 22770
rect 11870 22730 11880 22770
rect 11480 22720 11490 22730
rect 11400 22700 11490 22720
rect 11820 22710 11880 22730
rect 8740 22690 8800 22700
rect 7100 22640 7380 22680
rect 7420 22640 7430 22680
rect 7100 19490 7180 22640
rect 7370 22620 7430 22640
rect 7730 22670 8030 22680
rect 7730 22630 7880 22670
rect 7920 22630 7960 22670
rect 8000 22630 8030 22670
rect 7730 22620 8030 22630
rect 8140 22670 8320 22680
rect 8480 22670 8550 22690
rect 8140 22630 8260 22670
rect 8300 22630 8320 22670
rect 8140 22620 8320 22630
rect 8370 22630 8500 22670
rect 8540 22630 8550 22670
rect 8740 22670 8930 22690
rect 8740 22650 8800 22670
rect 8370 22610 8550 22630
rect 8730 22630 8800 22650
rect 8840 22630 8880 22670
rect 8920 22630 8930 22670
rect 8730 22610 8930 22630
rect 8970 22670 9070 22690
rect 8970 22630 9000 22670
rect 9040 22630 9070 22670
rect 8970 22610 9070 22630
rect 9200 22640 9220 22700
rect 9280 22640 9290 22700
rect 9200 22620 9290 22640
rect 9510 22670 9630 22690
rect 10560 22670 10620 22690
rect 11560 22670 11620 22690
rect 12710 22670 12950 22690
rect 9510 22630 9580 22670
rect 9620 22630 9630 22670
rect 9510 22610 9630 22630
rect 9930 22660 10230 22670
rect 9930 22620 10080 22660
rect 10120 22620 10160 22660
rect 10200 22620 10230 22660
rect 9930 22610 10230 22620
rect 10340 22660 10570 22670
rect 10340 22620 10460 22660
rect 10500 22630 10570 22660
rect 10610 22630 10620 22670
rect 10500 22620 10620 22630
rect 10340 22610 10620 22620
rect 10920 22660 11220 22670
rect 10920 22620 11070 22660
rect 11110 22620 11150 22660
rect 11190 22620 11220 22660
rect 10920 22610 11220 22620
rect 11330 22660 11570 22670
rect 11330 22620 11450 22660
rect 11490 22630 11570 22660
rect 11610 22630 11620 22670
rect 11490 22620 11620 22630
rect 11330 22610 11620 22620
rect 11920 22660 12220 22670
rect 11920 22620 12070 22660
rect 12110 22620 12150 22660
rect 12190 22620 12220 22660
rect 11920 22610 12220 22620
rect 12330 22660 12600 22670
rect 12330 22620 12450 22660
rect 12490 22620 12530 22660
rect 12570 22620 12600 22660
rect 12330 22610 12600 22620
rect 12710 22630 12820 22670
rect 12860 22630 12900 22670
rect 12940 22630 12950 22670
rect 12710 22610 12950 22630
rect 12990 22670 13180 22690
rect 12990 22630 13000 22670
rect 13040 22630 13130 22670
rect 13170 22630 13180 22670
rect 12990 22610 13180 22630
rect 13330 22670 13520 22690
rect 13330 22630 13340 22670
rect 13380 22630 13470 22670
rect 13510 22630 13520 22670
rect 13330 22610 13520 22630
rect 13890 22670 14080 22690
rect 13890 22630 13900 22670
rect 13940 22630 14030 22670
rect 14070 22630 14080 22670
rect 13890 22610 14080 22630
rect 14890 22670 15140 22690
rect 14890 22630 14900 22670
rect 14940 22630 15090 22670
rect 15130 22630 15140 22670
rect 14890 22610 15140 22630
rect 16830 22680 16960 22690
rect 16830 22630 16890 22680
rect 16940 22670 16960 22680
rect 17020 22670 17090 22690
rect 16940 22630 17040 22670
rect 17080 22630 17090 22670
rect 16830 22620 16960 22630
rect 17020 22610 17090 22630
rect 20540 22680 23140 22690
rect 20540 22630 20600 22680
rect 20650 22630 23140 22680
rect 20540 22620 23140 22630
rect 7460 22560 7540 22570
rect 7460 22520 7480 22560
rect 7520 22520 7540 22560
rect 7460 22510 7540 22520
rect 7720 22560 7800 22570
rect 7720 22520 7740 22560
rect 7780 22520 7800 22560
rect 7720 22510 7800 22520
rect 7480 21710 7520 22510
rect 7460 21700 7540 21710
rect 7460 21660 7480 21700
rect 7520 21660 7540 21700
rect 7740 21690 7780 22510
rect 7460 21650 7540 21660
rect 7720 21680 7800 21690
rect 7720 21640 7740 21680
rect 7780 21640 7800 21680
rect 7720 21630 7800 21640
rect 8370 21070 8420 22610
rect 8310 21010 8420 21070
rect 9510 21010 9550 22610
rect 13210 22570 13290 22580
rect 9660 22550 9740 22560
rect 9660 22510 9680 22550
rect 9720 22510 9740 22550
rect 9660 22500 9740 22510
rect 9920 22550 10000 22560
rect 9920 22510 9940 22550
rect 9980 22510 10000 22550
rect 9920 22500 10000 22510
rect 10650 22550 10730 22560
rect 10650 22510 10670 22550
rect 10710 22510 10730 22550
rect 10650 22500 10730 22510
rect 10910 22550 10990 22560
rect 10910 22510 10930 22550
rect 10970 22510 10990 22550
rect 10910 22500 10990 22510
rect 11650 22550 11730 22560
rect 11650 22510 11670 22550
rect 11710 22510 11730 22550
rect 11650 22500 11730 22510
rect 11910 22550 11990 22560
rect 11910 22510 11930 22550
rect 11970 22510 11990 22550
rect 13210 22530 13230 22570
rect 13270 22530 13290 22570
rect 13210 22520 13290 22530
rect 13550 22570 13630 22580
rect 13550 22530 13570 22570
rect 13610 22530 13630 22570
rect 13550 22520 13630 22530
rect 13770 22570 13850 22580
rect 13770 22530 13790 22570
rect 13830 22530 13850 22570
rect 13770 22520 13850 22530
rect 14110 22550 14190 22560
rect 11910 22500 11990 22510
rect 9680 21680 9720 22500
rect 9940 21680 9980 22500
rect 10670 21680 10710 22500
rect 10930 21680 10970 22500
rect 11670 21680 11710 22500
rect 11930 21680 11970 22500
rect 13230 21690 13270 22520
rect 13570 21690 13610 22520
rect 13790 21690 13830 22520
rect 14110 22510 14130 22550
rect 14170 22510 14190 22550
rect 14110 22500 14190 22510
rect 14330 22550 14410 22560
rect 14330 22510 14350 22550
rect 14390 22510 14410 22550
rect 14330 22500 14410 22510
rect 14550 22550 14630 22560
rect 14550 22510 14570 22550
rect 14610 22510 14630 22550
rect 14550 22500 14630 22510
rect 14770 22550 14850 22560
rect 14770 22510 14790 22550
rect 14830 22510 14850 22550
rect 14770 22500 14850 22510
rect 15170 22550 15250 22560
rect 15170 22510 15190 22550
rect 15230 22510 15250 22550
rect 15170 22500 15250 22510
rect 15390 22550 15470 22560
rect 15390 22510 15410 22550
rect 15450 22510 15470 22550
rect 15390 22500 15470 22510
rect 15610 22550 15690 22560
rect 15610 22510 15630 22550
rect 15670 22510 15690 22550
rect 15610 22500 15690 22510
rect 15830 22550 15910 22560
rect 15830 22510 15850 22550
rect 15890 22510 15910 22550
rect 15830 22500 15910 22510
rect 16050 22550 16130 22560
rect 16050 22510 16070 22550
rect 16110 22510 16130 22550
rect 16050 22500 16130 22510
rect 16270 22550 16350 22560
rect 16270 22510 16290 22550
rect 16330 22510 16350 22550
rect 16270 22500 16350 22510
rect 16490 22550 16570 22560
rect 16490 22510 16510 22550
rect 16550 22510 16570 22550
rect 16490 22500 16570 22510
rect 16710 22550 16790 22560
rect 16710 22510 16730 22550
rect 16770 22510 16790 22550
rect 16710 22500 16790 22510
rect 17120 22550 17200 22560
rect 17120 22510 17140 22550
rect 17180 22510 17200 22550
rect 17120 22500 17200 22510
rect 17340 22550 17420 22560
rect 17340 22510 17360 22550
rect 17400 22510 17420 22550
rect 17340 22500 17420 22510
rect 17560 22550 17640 22560
rect 17560 22510 17580 22550
rect 17620 22510 17640 22550
rect 17560 22500 17640 22510
rect 17780 22550 17860 22560
rect 17780 22510 17800 22550
rect 17840 22510 17860 22550
rect 17780 22500 17860 22510
rect 18000 22550 18080 22560
rect 18000 22510 18020 22550
rect 18060 22510 18080 22550
rect 18000 22500 18080 22510
rect 18220 22550 18300 22560
rect 18220 22510 18240 22550
rect 18280 22510 18300 22550
rect 18220 22500 18300 22510
rect 18440 22550 18520 22560
rect 18440 22510 18460 22550
rect 18500 22510 18520 22550
rect 18440 22500 18520 22510
rect 18660 22550 18740 22560
rect 18660 22510 18680 22550
rect 18720 22510 18740 22550
rect 18660 22500 18740 22510
rect 18880 22550 18960 22560
rect 18880 22510 18900 22550
rect 18940 22510 18960 22550
rect 18880 22500 18960 22510
rect 19100 22550 19180 22560
rect 19100 22510 19120 22550
rect 19160 22510 19180 22550
rect 19100 22500 19180 22510
rect 19320 22550 19400 22560
rect 19320 22510 19340 22550
rect 19380 22510 19400 22550
rect 19320 22500 19400 22510
rect 19540 22550 19620 22560
rect 19540 22510 19560 22550
rect 19600 22510 19620 22550
rect 19540 22500 19620 22510
rect 19760 22550 19840 22560
rect 19760 22510 19780 22550
rect 19820 22510 19840 22550
rect 19760 22500 19840 22510
rect 19980 22550 20060 22560
rect 19980 22510 20000 22550
rect 20040 22510 20060 22550
rect 19980 22500 20060 22510
rect 20200 22550 20280 22560
rect 20200 22510 20220 22550
rect 20260 22510 20280 22550
rect 20200 22500 20280 22510
rect 20420 22550 20500 22560
rect 20420 22510 20440 22550
rect 20480 22510 20500 22550
rect 20420 22500 20500 22510
rect 13210 21680 13290 21690
rect 9660 21670 9740 21680
rect 9660 21630 9680 21670
rect 9720 21630 9740 21670
rect 9660 21620 9740 21630
rect 9920 21670 10000 21680
rect 9920 21630 9940 21670
rect 9980 21630 10000 21670
rect 9920 21620 10000 21630
rect 10650 21670 10730 21680
rect 10650 21630 10670 21670
rect 10710 21630 10730 21670
rect 10650 21620 10730 21630
rect 10910 21670 10990 21680
rect 10910 21630 10930 21670
rect 10970 21630 10990 21670
rect 10910 21620 10990 21630
rect 11650 21670 11730 21680
rect 11650 21630 11670 21670
rect 11710 21630 11730 21670
rect 11650 21620 11730 21630
rect 11910 21670 11990 21680
rect 11910 21630 11930 21670
rect 11970 21630 11990 21670
rect 13210 21640 13230 21680
rect 13270 21640 13290 21680
rect 13210 21630 13290 21640
rect 13550 21680 13630 21690
rect 13550 21640 13570 21680
rect 13610 21640 13630 21680
rect 13550 21630 13630 21640
rect 13770 21680 13850 21690
rect 13770 21640 13790 21680
rect 13830 21640 13850 21680
rect 14130 21670 14170 22500
rect 14350 21670 14390 22500
rect 14570 21670 14610 22500
rect 14790 21670 14830 22500
rect 15190 21670 15230 22500
rect 15410 21670 15450 22500
rect 15630 21670 15670 22500
rect 15850 21670 15890 22500
rect 16070 21670 16110 22500
rect 16290 21670 16330 22500
rect 16510 21670 16550 22500
rect 16730 21670 16770 22500
rect 17140 21670 17180 22500
rect 17360 21670 17400 22500
rect 17580 21670 17620 22500
rect 17800 21670 17840 22500
rect 18020 21670 18060 22500
rect 18240 21670 18280 22500
rect 18460 21670 18500 22500
rect 18680 21670 18720 22500
rect 18900 21670 18940 22500
rect 19120 21670 19160 22500
rect 19340 21670 19380 22500
rect 19560 21670 19600 22500
rect 19780 21670 19820 22500
rect 20000 21670 20040 22500
rect 20220 21670 20260 22500
rect 20440 21670 20480 22500
rect 13770 21630 13850 21640
rect 14110 21660 14190 21670
rect 11910 21620 11990 21630
rect 14110 21620 14130 21660
rect 14170 21620 14190 21660
rect 14110 21610 14190 21620
rect 14330 21660 14410 21670
rect 14330 21620 14350 21660
rect 14390 21620 14410 21660
rect 14330 21610 14410 21620
rect 14550 21660 14630 21670
rect 14550 21620 14570 21660
rect 14610 21620 14630 21660
rect 14550 21610 14630 21620
rect 14770 21660 14850 21670
rect 14770 21620 14790 21660
rect 14830 21620 14850 21660
rect 14770 21610 14850 21620
rect 15170 21660 15250 21670
rect 15170 21620 15190 21660
rect 15230 21620 15250 21660
rect 15170 21610 15250 21620
rect 15390 21660 15470 21670
rect 15390 21620 15410 21660
rect 15450 21620 15470 21660
rect 15390 21610 15470 21620
rect 15610 21660 15690 21670
rect 15610 21620 15630 21660
rect 15670 21620 15690 21660
rect 15610 21610 15690 21620
rect 15830 21660 15910 21670
rect 15830 21620 15850 21660
rect 15890 21620 15910 21660
rect 15830 21610 15910 21620
rect 16050 21660 16130 21670
rect 16050 21620 16070 21660
rect 16110 21620 16130 21660
rect 16050 21610 16130 21620
rect 16270 21660 16350 21670
rect 16270 21620 16290 21660
rect 16330 21620 16350 21660
rect 16270 21610 16350 21620
rect 16490 21660 16570 21670
rect 16490 21620 16510 21660
rect 16550 21620 16570 21660
rect 16490 21610 16570 21620
rect 16710 21660 16790 21670
rect 16710 21620 16730 21660
rect 16770 21620 16790 21660
rect 16710 21610 16790 21620
rect 17120 21660 17200 21670
rect 17120 21620 17140 21660
rect 17180 21620 17200 21660
rect 17120 21610 17200 21620
rect 17340 21660 17420 21670
rect 17340 21620 17360 21660
rect 17400 21620 17420 21660
rect 17340 21610 17420 21620
rect 17560 21660 17640 21670
rect 17560 21620 17580 21660
rect 17620 21620 17640 21660
rect 17560 21610 17640 21620
rect 17780 21660 17860 21670
rect 17780 21620 17800 21660
rect 17840 21620 17860 21660
rect 17780 21610 17860 21620
rect 18000 21660 18080 21670
rect 18000 21620 18020 21660
rect 18060 21620 18080 21660
rect 18000 21610 18080 21620
rect 18220 21660 18300 21670
rect 18220 21620 18240 21660
rect 18280 21620 18300 21660
rect 18220 21610 18300 21620
rect 18440 21660 18520 21670
rect 18440 21620 18460 21660
rect 18500 21620 18520 21660
rect 18440 21610 18520 21620
rect 18660 21660 18740 21670
rect 18660 21620 18680 21660
rect 18720 21620 18740 21660
rect 18660 21610 18740 21620
rect 18880 21660 18960 21670
rect 18880 21620 18900 21660
rect 18940 21620 18960 21660
rect 18880 21610 18960 21620
rect 19100 21660 19180 21670
rect 19100 21620 19120 21660
rect 19160 21620 19180 21660
rect 19100 21610 19180 21620
rect 19320 21660 19400 21670
rect 19320 21620 19340 21660
rect 19380 21620 19400 21660
rect 19320 21610 19400 21620
rect 19540 21660 19620 21670
rect 19540 21620 19560 21660
rect 19600 21620 19620 21660
rect 19540 21610 19620 21620
rect 19760 21660 19840 21670
rect 19760 21620 19780 21660
rect 19820 21620 19840 21660
rect 19760 21610 19840 21620
rect 19980 21660 20060 21670
rect 19980 21620 20000 21660
rect 20040 21620 20060 21660
rect 19980 21610 20060 21620
rect 20200 21660 20280 21670
rect 20200 21620 20220 21660
rect 20260 21620 20280 21660
rect 20200 21610 20280 21620
rect 20420 21660 20500 21670
rect 20420 21620 20440 21660
rect 20480 21620 20500 21660
rect 20420 21610 20500 21620
rect 7280 21000 20640 21010
rect 7280 20960 7320 21000
rect 7360 20960 7400 21000
rect 7440 20960 7480 21000
rect 7520 20960 7560 21000
rect 7600 20960 7640 21000
rect 7680 20960 7720 21000
rect 7760 20960 7800 21000
rect 7840 20960 7880 21000
rect 7920 20960 7960 21000
rect 8000 20960 8040 21000
rect 8080 20960 8120 21000
rect 8160 20960 8200 21000
rect 8240 20960 8280 21000
rect 8320 20960 8360 21000
rect 8400 20960 8440 21000
rect 8480 20960 8520 21000
rect 8560 20960 8600 21000
rect 8640 20960 8680 21000
rect 8720 20960 8760 21000
rect 8800 20960 8840 21000
rect 8880 20960 8920 21000
rect 8960 20960 9000 21000
rect 9040 20960 9080 21000
rect 9120 20960 9160 21000
rect 9200 20960 9260 21000
rect 9300 20960 9340 21000
rect 9380 20960 9420 21000
rect 9460 20960 9500 21000
rect 9540 20960 9580 21000
rect 9620 20960 9660 21000
rect 9700 20960 9740 21000
rect 9780 20960 9820 21000
rect 9860 20960 9900 21000
rect 9940 20960 9980 21000
rect 10020 20960 10060 21000
rect 10100 20960 10140 21000
rect 10180 20960 10220 21000
rect 10260 20960 10300 21000
rect 10340 20960 10380 21000
rect 10420 20960 10460 21000
rect 10500 20960 10540 21000
rect 10580 20960 10620 21000
rect 10660 20960 10700 21000
rect 10740 20960 10780 21000
rect 10820 20960 10860 21000
rect 10900 20960 10940 21000
rect 10980 20960 11020 21000
rect 11060 20960 11100 21000
rect 11140 20960 11180 21000
rect 11220 20960 11260 21000
rect 11300 20960 11340 21000
rect 11380 20960 11420 21000
rect 11460 20960 11500 21000
rect 11540 20960 11580 21000
rect 11620 20960 11660 21000
rect 11700 20960 11740 21000
rect 11780 20960 11820 21000
rect 11860 20960 11900 21000
rect 11940 20960 11980 21000
rect 12020 20960 12060 21000
rect 12100 20960 12140 21000
rect 12180 20960 12220 21000
rect 12260 20960 12300 21000
rect 12340 20960 12380 21000
rect 12420 20960 12460 21000
rect 12500 20960 12540 21000
rect 12580 20960 12620 21000
rect 12660 20960 12700 21000
rect 12740 20960 12780 21000
rect 12820 20960 12880 21000
rect 12920 20960 12960 21000
rect 13000 20960 13040 21000
rect 13080 20960 13120 21000
rect 13160 20960 13200 21000
rect 13240 20960 13280 21000
rect 13320 20960 13360 21000
rect 13400 20960 13440 21000
rect 13480 20960 13520 21000
rect 13560 20960 13600 21000
rect 13640 20960 13680 21000
rect 13720 20960 13760 21000
rect 13800 20960 13840 21000
rect 13880 20960 13920 21000
rect 13960 20960 14000 21000
rect 14040 20960 14080 21000
rect 14120 20960 14160 21000
rect 14200 20960 14240 21000
rect 14280 20960 14320 21000
rect 14360 20960 14400 21000
rect 14440 20960 14480 21000
rect 14520 20960 14560 21000
rect 14600 20960 14640 21000
rect 14680 20960 14720 21000
rect 14760 20960 14800 21000
rect 14840 20960 14880 21000
rect 14920 20960 14960 21000
rect 15000 20960 15040 21000
rect 15080 20960 15120 21000
rect 15160 20960 15200 21000
rect 15240 20960 15280 21000
rect 15320 20960 15360 21000
rect 15400 20960 15440 21000
rect 15480 20960 15520 21000
rect 15560 20960 15600 21000
rect 15640 20960 15680 21000
rect 15720 20960 15760 21000
rect 15800 20960 15840 21000
rect 15880 20960 15920 21000
rect 15960 20960 16000 21000
rect 16040 20960 16080 21000
rect 16120 20960 16160 21000
rect 16200 20960 16240 21000
rect 16280 20960 16320 21000
rect 16360 20960 16400 21000
rect 16440 20960 16480 21000
rect 16520 20960 16560 21000
rect 16600 20960 16640 21000
rect 16680 20960 16720 21000
rect 16760 20960 16800 21000
rect 16840 20960 16880 21000
rect 16920 20960 16960 21000
rect 17000 20960 17040 21000
rect 17080 20960 17120 21000
rect 17160 20960 17200 21000
rect 17240 20960 17280 21000
rect 17320 20960 17360 21000
rect 17400 20960 17440 21000
rect 17480 20960 17520 21000
rect 17560 20960 17600 21000
rect 17640 20960 17680 21000
rect 17720 20960 17760 21000
rect 17800 20960 17840 21000
rect 17880 20960 17920 21000
rect 17960 20960 18000 21000
rect 18040 20960 18080 21000
rect 18120 20960 18160 21000
rect 18200 20960 18240 21000
rect 18280 20960 18320 21000
rect 18360 20960 18400 21000
rect 18440 20960 18480 21000
rect 18520 20960 18560 21000
rect 18600 20960 18640 21000
rect 18680 20960 18720 21000
rect 18760 20960 18800 21000
rect 18840 20960 18880 21000
rect 18920 20960 18960 21000
rect 19000 20960 19040 21000
rect 19080 20960 19120 21000
rect 19160 20960 19200 21000
rect 19240 20960 19280 21000
rect 19320 20960 19360 21000
rect 19400 20960 19440 21000
rect 19480 20960 19520 21000
rect 19560 20960 19600 21000
rect 19640 20960 19680 21000
rect 19720 20960 19760 21000
rect 19800 20960 19840 21000
rect 19880 20960 19920 21000
rect 19960 20960 20000 21000
rect 20040 20960 20080 21000
rect 20120 20960 20160 21000
rect 20200 20960 20240 21000
rect 20280 20960 20320 21000
rect 20360 20960 20400 21000
rect 20440 20960 20480 21000
rect 20520 20960 20560 21000
rect 20600 20960 20640 21000
rect 7280 20890 20640 20960
rect 7280 20480 17670 20890
rect 7280 20470 8230 20480
rect 7280 20430 7320 20470
rect 7360 20430 7400 20470
rect 7440 20430 7480 20470
rect 7520 20430 7560 20470
rect 7600 20430 7640 20470
rect 7680 20430 7720 20470
rect 7760 20430 7800 20470
rect 7840 20430 7880 20470
rect 7920 20430 7960 20470
rect 8000 20430 8040 20470
rect 8080 20430 8120 20470
rect 8160 20430 8230 20470
rect 7280 20420 8230 20430
rect 8360 20410 17670 20480
rect 8360 20350 12730 20410
rect 12800 20350 17670 20410
rect 8360 20090 17670 20350
rect 18500 20090 20640 20890
rect 8360 20030 20640 20090
rect 8310 20020 20640 20030
rect 8310 19980 8360 20020
rect 8400 19980 8440 20020
rect 8480 19980 8520 20020
rect 8560 19980 8600 20020
rect 8640 19980 8680 20020
rect 8720 19980 8760 20020
rect 8800 19980 8840 20020
rect 8880 19980 8920 20020
rect 8960 19980 9000 20020
rect 9040 19980 9080 20020
rect 9120 19980 9160 20020
rect 9200 19980 9260 20020
rect 9300 19980 9340 20020
rect 9380 19980 9420 20020
rect 9460 19980 9500 20020
rect 9540 19980 9580 20020
rect 9620 19980 9660 20020
rect 9700 19980 9740 20020
rect 9780 19980 9820 20020
rect 9860 19980 9900 20020
rect 9940 19980 9980 20020
rect 10020 19980 10060 20020
rect 10100 19980 10140 20020
rect 10180 19980 10220 20020
rect 10260 19980 10300 20020
rect 10340 19980 10380 20020
rect 10420 19980 10460 20020
rect 10500 19980 10540 20020
rect 10580 19980 10620 20020
rect 10660 19980 10700 20020
rect 10740 19980 10780 20020
rect 10820 19980 10860 20020
rect 10900 19980 10940 20020
rect 10980 19980 11020 20020
rect 11060 19980 11100 20020
rect 11140 19980 11180 20020
rect 11220 19980 11260 20020
rect 11300 19980 11340 20020
rect 11380 19980 11420 20020
rect 11460 19980 11500 20020
rect 11540 19980 11580 20020
rect 11620 19980 11660 20020
rect 11700 19980 11740 20020
rect 11780 19980 11820 20020
rect 11860 19980 11900 20020
rect 11940 19980 11980 20020
rect 12020 19980 12060 20020
rect 12100 19980 12140 20020
rect 12180 19980 12220 20020
rect 12260 19980 12300 20020
rect 12340 19980 12380 20020
rect 12420 19980 12460 20020
rect 12500 19980 12540 20020
rect 12580 19980 12620 20020
rect 12660 19980 12700 20020
rect 12740 19980 12780 20020
rect 12820 19980 12860 20020
rect 12900 19980 12940 20020
rect 12980 19980 13040 20020
rect 13080 19980 13120 20020
rect 13160 19980 13200 20020
rect 13240 19980 13280 20020
rect 13320 19980 13360 20020
rect 13400 19980 13440 20020
rect 13480 19980 13520 20020
rect 13560 19980 13600 20020
rect 13640 19980 13680 20020
rect 13720 19980 13760 20020
rect 13800 19980 13840 20020
rect 13880 19980 13920 20020
rect 13960 19980 14000 20020
rect 14040 19980 14080 20020
rect 14120 19980 14160 20020
rect 14200 19980 14240 20020
rect 14280 19980 14320 20020
rect 14360 19980 14400 20020
rect 14440 19980 14480 20020
rect 14520 19980 14560 20020
rect 14600 19980 14640 20020
rect 14680 19980 14720 20020
rect 14760 19980 14800 20020
rect 14840 19980 14880 20020
rect 14920 19980 14960 20020
rect 15000 19980 15040 20020
rect 15080 19980 15120 20020
rect 15160 19980 15200 20020
rect 15240 19980 15280 20020
rect 15320 19980 15360 20020
rect 15400 19980 15440 20020
rect 15480 19980 15520 20020
rect 15560 19980 15600 20020
rect 15640 19980 15680 20020
rect 15720 19980 15760 20020
rect 15800 19980 15840 20020
rect 15880 19980 15920 20020
rect 15960 19980 16000 20020
rect 16040 19980 16080 20020
rect 16120 19980 16160 20020
rect 16200 19980 16240 20020
rect 16280 19980 16320 20020
rect 16360 19980 16400 20020
rect 16440 19980 16480 20020
rect 16520 19980 16560 20020
rect 16600 19980 16640 20020
rect 16680 19980 16720 20020
rect 16760 19980 16800 20020
rect 16840 19980 16880 20020
rect 16920 19980 16960 20020
rect 17000 19980 17040 20020
rect 17080 19980 17120 20020
rect 17160 19980 17200 20020
rect 17240 19980 17280 20020
rect 17320 19980 17360 20020
rect 17400 19980 17440 20020
rect 17480 19980 17520 20020
rect 17560 19980 17600 20020
rect 17640 19980 17680 20020
rect 17720 19980 17760 20020
rect 17800 19980 17840 20020
rect 17880 19980 17920 20020
rect 17960 19980 18000 20020
rect 18040 19980 18080 20020
rect 18120 19980 18160 20020
rect 18200 19980 18240 20020
rect 18280 19980 18320 20020
rect 18360 19980 18400 20020
rect 18440 19980 18480 20020
rect 18520 19980 18560 20020
rect 18600 19980 18640 20020
rect 18680 19980 18720 20020
rect 18760 19980 18800 20020
rect 18840 19980 18880 20020
rect 18920 19980 18960 20020
rect 19000 19980 19040 20020
rect 19080 19980 19120 20020
rect 19160 19980 19200 20020
rect 19240 19980 19280 20020
rect 19320 19980 19360 20020
rect 19400 19980 19440 20020
rect 19480 19980 19520 20020
rect 19560 19980 19600 20020
rect 19640 19980 19680 20020
rect 19720 19980 19760 20020
rect 19800 19980 19840 20020
rect 19880 19980 19920 20020
rect 19960 19980 20000 20020
rect 20040 19980 20080 20020
rect 20120 19980 20160 20020
rect 20200 19980 20240 20020
rect 20280 19980 20320 20020
rect 20360 19980 20400 20020
rect 20440 19980 20480 20020
rect 20520 19980 20560 20020
rect 20600 19980 20640 20020
rect 8310 19970 20640 19980
rect 8310 19910 8420 19970
rect 7090 19470 7190 19490
rect 7090 19410 7110 19470
rect 7170 19410 7190 19470
rect 7090 19390 7190 19410
rect 6940 18620 6960 18680
rect 7020 18620 7040 18680
rect 6940 18600 7040 18620
rect 7100 18190 7180 19390
rect 7350 19310 7490 19320
rect 7350 19270 7400 19310
rect 7440 19270 7490 19310
rect 7350 19260 7490 19270
rect 7400 18440 7440 19260
rect 7210 18420 7310 18440
rect 7210 18360 7230 18420
rect 7290 18360 7310 18420
rect 7350 18430 7490 18440
rect 7350 18390 7400 18430
rect 7440 18390 7490 18430
rect 7350 18380 7490 18390
rect 7210 18340 7310 18360
rect 8370 18370 8420 19910
rect 9660 19360 9740 19370
rect 9660 19320 9680 19360
rect 9720 19320 9740 19360
rect 9660 19310 9740 19320
rect 9920 19360 10000 19370
rect 9920 19320 9940 19360
rect 9980 19320 10000 19360
rect 9920 19310 10000 19320
rect 10650 19360 10730 19370
rect 10650 19320 10670 19360
rect 10710 19320 10730 19360
rect 10650 19310 10730 19320
rect 10910 19360 10990 19370
rect 10910 19320 10930 19360
rect 10970 19320 10990 19360
rect 10910 19310 10990 19320
rect 11650 19350 11730 19360
rect 11650 19310 11670 19350
rect 11710 19310 11730 19350
rect 9680 18480 9720 19310
rect 9940 18480 9980 19310
rect 10670 18480 10710 19310
rect 10930 18480 10970 19310
rect 11650 19300 11730 19310
rect 9660 18470 9740 18480
rect 9660 18430 9680 18470
rect 9720 18430 9740 18470
rect 9660 18420 9740 18430
rect 9920 18470 10000 18480
rect 9920 18430 9940 18470
rect 9980 18430 10000 18470
rect 9920 18420 10000 18430
rect 10650 18470 10730 18480
rect 10650 18430 10670 18470
rect 10710 18430 10730 18470
rect 10650 18420 10730 18430
rect 10910 18470 10990 18480
rect 11670 18470 11710 19300
rect 10910 18430 10930 18470
rect 10970 18430 10990 18470
rect 10910 18420 10990 18430
rect 11650 18460 11730 18470
rect 11650 18420 11670 18460
rect 11710 18420 11730 18460
rect 11650 18410 11730 18420
rect 8370 18350 8550 18370
rect 7230 18300 7290 18340
rect 8370 18310 8500 18350
rect 8540 18310 8550 18350
rect 8730 18350 8930 18370
rect 8730 18330 8800 18350
rect 7230 18280 7610 18300
rect 7230 18240 7560 18280
rect 7600 18240 7610 18280
rect 7230 18220 7610 18240
rect 7890 18280 8020 18300
rect 8480 18290 8550 18310
rect 8740 18310 8800 18330
rect 8840 18310 8880 18350
rect 8920 18310 8930 18350
rect 8740 18290 8930 18310
rect 8970 18350 9070 18370
rect 9470 18350 9630 18370
rect 8970 18310 9000 18350
rect 9040 18310 9070 18350
rect 8970 18290 9070 18310
rect 9200 18330 9290 18350
rect 7890 18240 7970 18280
rect 8010 18240 8020 18280
rect 8630 18270 8700 18290
rect 8740 18280 8800 18290
rect 8630 18260 8650 18270
rect 7890 18220 8020 18240
rect 8360 18230 8650 18260
rect 8690 18230 8700 18270
rect 9200 18270 9220 18330
rect 9280 18270 9290 18330
rect 9200 18250 9290 18270
rect 9470 18310 9580 18350
rect 9620 18310 9630 18350
rect 9930 18360 10230 18370
rect 9930 18320 10080 18360
rect 10120 18320 10160 18360
rect 10200 18320 10230 18360
rect 9930 18310 10230 18320
rect 10340 18360 10620 18370
rect 10340 18320 10460 18360
rect 10500 18350 10620 18360
rect 10500 18320 10570 18350
rect 10340 18310 10570 18320
rect 10610 18310 10620 18350
rect 10920 18360 11220 18370
rect 10920 18320 11070 18360
rect 11110 18320 11150 18360
rect 11190 18320 11220 18360
rect 10920 18310 11220 18320
rect 11330 18360 11620 18370
rect 11330 18320 11450 18360
rect 11490 18350 11620 18360
rect 11490 18320 11570 18350
rect 11330 18310 11570 18320
rect 11610 18310 11620 18350
rect 9470 18290 9630 18310
rect 10560 18290 10620 18310
rect 11560 18290 11620 18310
rect 7100 18170 7350 18190
rect 7100 18130 7300 18170
rect 7340 18130 7350 18170
rect 7100 18110 7350 18130
rect 7890 18080 7950 18220
rect 8360 18210 8700 18230
rect 8360 18080 8410 18210
rect 9080 18180 9170 18200
rect 9080 18130 9100 18180
rect 9150 18130 9170 18180
rect 9080 18110 9170 18130
rect 9470 18120 9540 18290
rect 9830 18250 9890 18270
rect 9830 18210 9840 18250
rect 9880 18210 9890 18250
rect 9830 18190 9890 18210
rect 10400 18260 10490 18280
rect 11770 18270 11820 19970
rect 14110 19360 14190 19370
rect 11910 19350 11990 19360
rect 11910 19310 11930 19350
rect 11970 19310 11990 19350
rect 11910 19300 11990 19310
rect 13210 19340 13290 19350
rect 13210 19300 13230 19340
rect 13270 19300 13290 19340
rect 11930 18470 11970 19300
rect 13210 19290 13290 19300
rect 13550 19340 13630 19350
rect 13550 19300 13570 19340
rect 13610 19300 13630 19340
rect 13550 19290 13630 19300
rect 13770 19340 13850 19350
rect 13770 19300 13790 19340
rect 13830 19300 13850 19340
rect 14110 19320 14130 19360
rect 14170 19320 14190 19360
rect 14110 19310 14190 19320
rect 14330 19360 14410 19370
rect 14330 19320 14350 19360
rect 14390 19320 14410 19360
rect 14330 19310 14410 19320
rect 14550 19360 14630 19370
rect 14550 19320 14570 19360
rect 14610 19320 14630 19360
rect 14550 19310 14630 19320
rect 14770 19360 14850 19370
rect 14770 19320 14790 19360
rect 14830 19320 14850 19360
rect 14770 19310 14850 19320
rect 15170 19360 15250 19370
rect 15170 19320 15190 19360
rect 15230 19320 15250 19360
rect 15170 19310 15250 19320
rect 15390 19360 15470 19370
rect 15390 19320 15410 19360
rect 15450 19320 15470 19360
rect 15390 19310 15470 19320
rect 15610 19360 15690 19370
rect 15610 19320 15630 19360
rect 15670 19320 15690 19360
rect 15610 19310 15690 19320
rect 15830 19360 15910 19370
rect 15830 19320 15850 19360
rect 15890 19320 15910 19360
rect 15830 19310 15910 19320
rect 16050 19360 16130 19370
rect 16050 19320 16070 19360
rect 16110 19320 16130 19360
rect 16050 19310 16130 19320
rect 16270 19360 16350 19370
rect 16270 19320 16290 19360
rect 16330 19320 16350 19360
rect 16270 19310 16350 19320
rect 16490 19360 16570 19370
rect 16490 19320 16510 19360
rect 16550 19320 16570 19360
rect 16490 19310 16570 19320
rect 16710 19360 16790 19370
rect 16710 19320 16730 19360
rect 16770 19320 16790 19360
rect 16710 19310 16790 19320
rect 17120 19360 17200 19370
rect 17120 19320 17140 19360
rect 17180 19320 17200 19360
rect 17120 19310 17200 19320
rect 17340 19360 17420 19370
rect 17340 19320 17360 19360
rect 17400 19320 17420 19360
rect 17340 19310 17420 19320
rect 17560 19360 17640 19370
rect 17560 19320 17580 19360
rect 17620 19320 17640 19360
rect 17560 19310 17640 19320
rect 17780 19360 17860 19370
rect 17780 19320 17800 19360
rect 17840 19320 17860 19360
rect 17780 19310 17860 19320
rect 18000 19360 18080 19370
rect 18000 19320 18020 19360
rect 18060 19320 18080 19360
rect 18000 19310 18080 19320
rect 18220 19360 18300 19370
rect 18220 19320 18240 19360
rect 18280 19320 18300 19360
rect 18220 19310 18300 19320
rect 18440 19360 18520 19370
rect 18440 19320 18460 19360
rect 18500 19320 18520 19360
rect 18440 19310 18520 19320
rect 18660 19360 18740 19370
rect 18660 19320 18680 19360
rect 18720 19320 18740 19360
rect 18660 19310 18740 19320
rect 18880 19360 18960 19370
rect 18880 19320 18900 19360
rect 18940 19320 18960 19360
rect 18880 19310 18960 19320
rect 19100 19360 19180 19370
rect 19100 19320 19120 19360
rect 19160 19320 19180 19360
rect 19100 19310 19180 19320
rect 19320 19360 19400 19370
rect 19320 19320 19340 19360
rect 19380 19320 19400 19360
rect 19320 19310 19400 19320
rect 19540 19360 19620 19370
rect 19540 19320 19560 19360
rect 19600 19320 19620 19360
rect 19540 19310 19620 19320
rect 19760 19360 19840 19370
rect 19760 19320 19780 19360
rect 19820 19320 19840 19360
rect 19760 19310 19840 19320
rect 19980 19360 20060 19370
rect 19980 19320 20000 19360
rect 20040 19320 20060 19360
rect 19980 19310 20060 19320
rect 20200 19360 20280 19370
rect 20200 19320 20220 19360
rect 20260 19320 20280 19360
rect 20200 19310 20280 19320
rect 20420 19360 20500 19370
rect 20420 19320 20440 19360
rect 20480 19320 20500 19360
rect 20420 19310 20500 19320
rect 13770 19290 13850 19300
rect 11910 18460 11990 18470
rect 13230 18460 13270 19290
rect 13570 18460 13610 19290
rect 13790 18460 13830 19290
rect 14130 18480 14170 19310
rect 14350 18480 14390 19310
rect 14570 18480 14610 19310
rect 14790 18480 14830 19310
rect 15190 18480 15230 19310
rect 15410 18480 15450 19310
rect 15630 18480 15670 19310
rect 15850 18480 15890 19310
rect 16070 18480 16110 19310
rect 16290 18480 16330 19310
rect 16510 18480 16550 19310
rect 16730 18480 16770 19310
rect 17140 18480 17180 19310
rect 17360 18480 17400 19310
rect 17580 18480 17620 19310
rect 17800 18480 17840 19310
rect 18020 18480 18060 19310
rect 18240 18480 18280 19310
rect 18460 18480 18500 19310
rect 18680 18480 18720 19310
rect 18900 18480 18940 19310
rect 19120 18480 19160 19310
rect 19340 18480 19380 19310
rect 19560 18480 19600 19310
rect 19780 18480 19820 19310
rect 20000 18480 20040 19310
rect 20220 18480 20260 19310
rect 20440 18480 20480 19310
rect 14110 18470 14190 18480
rect 11910 18420 11930 18460
rect 11970 18420 11990 18460
rect 11910 18410 11990 18420
rect 13210 18450 13290 18460
rect 13210 18410 13230 18450
rect 13270 18410 13290 18450
rect 13210 18400 13290 18410
rect 13550 18450 13630 18460
rect 13550 18410 13570 18450
rect 13610 18410 13630 18450
rect 13550 18400 13630 18410
rect 13770 18450 13850 18460
rect 13770 18410 13790 18450
rect 13830 18410 13850 18450
rect 14110 18430 14130 18470
rect 14170 18430 14190 18470
rect 14110 18420 14190 18430
rect 14330 18470 14410 18480
rect 14330 18430 14350 18470
rect 14390 18430 14410 18470
rect 14330 18420 14410 18430
rect 14550 18470 14630 18480
rect 14550 18430 14570 18470
rect 14610 18430 14630 18470
rect 14550 18420 14630 18430
rect 14770 18470 14850 18480
rect 14770 18430 14790 18470
rect 14830 18430 14850 18470
rect 14770 18420 14850 18430
rect 15170 18470 15250 18480
rect 15170 18430 15190 18470
rect 15230 18430 15250 18470
rect 15170 18420 15250 18430
rect 15390 18470 15470 18480
rect 15390 18430 15410 18470
rect 15450 18430 15470 18470
rect 15390 18420 15470 18430
rect 15610 18470 15690 18480
rect 15610 18430 15630 18470
rect 15670 18430 15690 18470
rect 15610 18420 15690 18430
rect 15830 18470 15910 18480
rect 15830 18430 15850 18470
rect 15890 18430 15910 18470
rect 15830 18420 15910 18430
rect 16050 18470 16130 18480
rect 16050 18430 16070 18470
rect 16110 18430 16130 18470
rect 16050 18420 16130 18430
rect 16270 18470 16350 18480
rect 16270 18430 16290 18470
rect 16330 18430 16350 18470
rect 16270 18420 16350 18430
rect 16490 18470 16570 18480
rect 16490 18430 16510 18470
rect 16550 18430 16570 18470
rect 16490 18420 16570 18430
rect 16710 18470 16790 18480
rect 16710 18430 16730 18470
rect 16770 18430 16790 18470
rect 16710 18420 16790 18430
rect 17120 18470 17200 18480
rect 17120 18430 17140 18470
rect 17180 18430 17200 18470
rect 17120 18420 17200 18430
rect 17340 18470 17420 18480
rect 17340 18430 17360 18470
rect 17400 18430 17420 18470
rect 17340 18420 17420 18430
rect 17560 18470 17640 18480
rect 17560 18430 17580 18470
rect 17620 18430 17640 18470
rect 17560 18420 17640 18430
rect 17780 18470 17860 18480
rect 17780 18430 17800 18470
rect 17840 18430 17860 18470
rect 17780 18420 17860 18430
rect 18000 18470 18080 18480
rect 18000 18430 18020 18470
rect 18060 18430 18080 18470
rect 18000 18420 18080 18430
rect 18220 18470 18300 18480
rect 18220 18430 18240 18470
rect 18280 18430 18300 18470
rect 18220 18420 18300 18430
rect 18440 18470 18520 18480
rect 18440 18430 18460 18470
rect 18500 18430 18520 18470
rect 18440 18420 18520 18430
rect 18660 18470 18740 18480
rect 18660 18430 18680 18470
rect 18720 18430 18740 18470
rect 18660 18420 18740 18430
rect 18880 18470 18960 18480
rect 18880 18430 18900 18470
rect 18940 18430 18960 18470
rect 18880 18420 18960 18430
rect 19100 18470 19180 18480
rect 19100 18430 19120 18470
rect 19160 18430 19180 18470
rect 19100 18420 19180 18430
rect 19320 18470 19400 18480
rect 19320 18430 19340 18470
rect 19380 18430 19400 18470
rect 19320 18420 19400 18430
rect 19540 18470 19620 18480
rect 19540 18430 19560 18470
rect 19600 18430 19620 18470
rect 19540 18420 19620 18430
rect 19760 18470 19840 18480
rect 19760 18430 19780 18470
rect 19820 18430 19840 18470
rect 19760 18420 19840 18430
rect 19980 18470 20060 18480
rect 19980 18430 20000 18470
rect 20040 18430 20060 18470
rect 19980 18420 20060 18430
rect 20200 18470 20280 18480
rect 20200 18430 20220 18470
rect 20260 18430 20280 18470
rect 20200 18420 20280 18430
rect 20420 18470 20500 18480
rect 20420 18430 20440 18470
rect 20480 18430 20500 18470
rect 20420 18420 20500 18430
rect 13770 18400 13850 18410
rect 11920 18360 12220 18370
rect 11920 18320 12070 18360
rect 12110 18320 12150 18360
rect 12190 18320 12220 18360
rect 11920 18310 12220 18320
rect 12330 18360 12600 18370
rect 12330 18320 12450 18360
rect 12490 18320 12530 18360
rect 12570 18320 12600 18360
rect 12330 18310 12600 18320
rect 12710 18350 12950 18370
rect 12710 18310 12820 18350
rect 12860 18310 12900 18350
rect 12940 18310 12950 18350
rect 12710 18290 12950 18310
rect 12990 18350 13180 18370
rect 12990 18310 13000 18350
rect 13040 18310 13130 18350
rect 13170 18310 13180 18350
rect 12990 18290 13180 18310
rect 13330 18350 13520 18370
rect 13330 18310 13340 18350
rect 13380 18310 13470 18350
rect 13510 18310 13520 18350
rect 13330 18290 13520 18310
rect 13890 18350 14080 18370
rect 13890 18310 13900 18350
rect 13940 18310 14030 18350
rect 14070 18310 14080 18350
rect 13890 18290 14080 18310
rect 14890 18350 15140 18370
rect 14890 18310 14900 18350
rect 14940 18310 15090 18350
rect 15130 18310 15140 18350
rect 14890 18290 15140 18310
rect 16830 18350 16960 18360
rect 17020 18350 17090 18370
rect 16830 18300 16890 18350
rect 16940 18310 17040 18350
rect 17080 18310 17090 18350
rect 16940 18300 16960 18310
rect 16830 18290 16960 18300
rect 17020 18290 17090 18310
rect 20540 18350 22860 18360
rect 20540 18300 20600 18350
rect 20650 18300 22860 18350
rect 20540 18290 22860 18300
rect 10400 18200 10410 18260
rect 10480 18250 10490 18260
rect 10820 18250 10880 18270
rect 10480 18210 10830 18250
rect 10870 18210 10880 18250
rect 10480 18200 10490 18210
rect 10400 18180 10490 18200
rect 10820 18190 10880 18210
rect 11770 18250 11880 18270
rect 11770 18210 11830 18250
rect 11870 18210 11880 18250
rect 11770 18200 11880 18210
rect 11820 18190 11880 18200
rect 7760 18070 7950 18080
rect 7760 18030 7780 18070
rect 7820 18030 7950 18070
rect 7760 18020 7950 18030
rect 8120 18070 8410 18080
rect 8120 18030 8190 18070
rect 8230 18030 8410 18070
rect 8120 18020 8410 18030
rect 9090 17980 9160 18110
rect 9460 18100 9550 18120
rect 9460 18040 9470 18100
rect 9540 18040 9550 18100
rect 9460 18020 9550 18040
rect 9080 17960 9170 17980
rect 9080 17900 9090 17960
rect 9160 17900 9170 17960
rect 9080 17880 9170 17900
rect 7280 17700 20620 17710
rect 7280 17660 7320 17700
rect 7360 17660 7400 17700
rect 7440 17660 7480 17700
rect 7520 17660 7560 17700
rect 7600 17660 7640 17700
rect 7680 17660 7720 17700
rect 7760 17660 7800 17700
rect 7840 17660 7880 17700
rect 7920 17660 7960 17700
rect 8000 17660 8040 17700
rect 8080 17660 8120 17700
rect 8160 17660 8200 17700
rect 8240 17660 8280 17700
rect 8320 17660 8360 17700
rect 8400 17660 8440 17700
rect 8480 17660 8520 17700
rect 8560 17660 8600 17700
rect 8640 17660 8680 17700
rect 8720 17660 8760 17700
rect 8800 17660 8840 17700
rect 8880 17660 8920 17700
rect 8960 17660 9000 17700
rect 9040 17660 9080 17700
rect 9120 17660 9160 17700
rect 9200 17660 9270 17700
rect 9310 17660 9350 17700
rect 9390 17660 9430 17700
rect 9470 17660 9510 17700
rect 9550 17660 9590 17700
rect 9630 17660 9670 17700
rect 9710 17660 9750 17700
rect 9790 17660 9830 17700
rect 9870 17660 9910 17700
rect 9950 17660 9990 17700
rect 10030 17660 10070 17700
rect 10110 17660 10150 17700
rect 10190 17660 10230 17700
rect 10270 17660 10310 17700
rect 10350 17660 10390 17700
rect 10430 17660 10470 17700
rect 10510 17660 10550 17700
rect 10590 17660 10630 17700
rect 10670 17660 10710 17700
rect 10750 17660 10790 17700
rect 10830 17660 10870 17700
rect 10910 17660 10950 17700
rect 10990 17660 11030 17700
rect 11070 17660 11110 17700
rect 11150 17660 11190 17700
rect 11230 17660 11270 17700
rect 11310 17660 11350 17700
rect 11390 17660 11430 17700
rect 11470 17660 11510 17700
rect 11550 17660 11590 17700
rect 11630 17660 11670 17700
rect 11710 17660 11750 17700
rect 11790 17660 11830 17700
rect 11870 17660 11910 17700
rect 11950 17660 11990 17700
rect 12030 17660 12070 17700
rect 12110 17660 12150 17700
rect 12190 17660 12230 17700
rect 12270 17660 12310 17700
rect 12350 17660 12390 17700
rect 12430 17660 12470 17700
rect 12510 17660 12550 17700
rect 12590 17660 12630 17700
rect 12670 17660 12710 17700
rect 12750 17660 12790 17700
rect 12830 17660 12870 17700
rect 12910 17660 12950 17700
rect 12990 17660 13030 17700
rect 13070 17660 13110 17700
rect 13150 17660 13190 17700
rect 13230 17660 13270 17700
rect 13310 17660 13350 17700
rect 13390 17660 13430 17700
rect 13470 17660 13510 17700
rect 13550 17660 13590 17700
rect 13630 17660 13670 17700
rect 13710 17660 13750 17700
rect 13790 17660 13830 17700
rect 13870 17660 13910 17700
rect 13950 17660 13990 17700
rect 14030 17660 14070 17700
rect 14110 17660 14150 17700
rect 14190 17660 14230 17700
rect 14270 17660 14310 17700
rect 14350 17660 14390 17700
rect 14430 17660 14470 17700
rect 14510 17660 14550 17700
rect 14590 17660 14630 17700
rect 14670 17660 14710 17700
rect 14750 17660 14790 17700
rect 14830 17660 14870 17700
rect 14910 17660 14950 17700
rect 14990 17660 15030 17700
rect 15070 17660 15110 17700
rect 15150 17660 15190 17700
rect 15230 17660 15270 17700
rect 15310 17660 15350 17700
rect 15390 17660 15430 17700
rect 15470 17660 15510 17700
rect 15550 17660 15590 17700
rect 15630 17660 15670 17700
rect 15710 17660 15750 17700
rect 15790 17660 15830 17700
rect 15870 17660 15910 17700
rect 15950 17660 15990 17700
rect 16030 17660 16070 17700
rect 16110 17660 16150 17700
rect 16190 17660 16230 17700
rect 16270 17660 16310 17700
rect 16350 17660 16390 17700
rect 16430 17660 16470 17700
rect 16510 17660 16550 17700
rect 16590 17660 16630 17700
rect 16670 17660 16710 17700
rect 16750 17660 16790 17700
rect 16830 17660 16870 17700
rect 16910 17660 16950 17700
rect 16990 17660 17030 17700
rect 17070 17660 17110 17700
rect 17150 17660 17190 17700
rect 17230 17660 17270 17700
rect 17310 17660 17350 17700
rect 17390 17660 17430 17700
rect 17470 17660 17510 17700
rect 17550 17660 17590 17700
rect 17630 17660 17670 17700
rect 17710 17660 17750 17700
rect 17790 17660 17830 17700
rect 17870 17660 17910 17700
rect 17950 17660 17990 17700
rect 18030 17660 18070 17700
rect 18110 17660 18150 17700
rect 18190 17660 18230 17700
rect 18270 17660 18310 17700
rect 18350 17660 18390 17700
rect 18430 17660 18470 17700
rect 18510 17660 18550 17700
rect 18590 17660 18630 17700
rect 18670 17660 18710 17700
rect 18750 17660 18790 17700
rect 18830 17660 18870 17700
rect 18910 17660 18950 17700
rect 18990 17660 19030 17700
rect 19070 17660 19110 17700
rect 19150 17660 19190 17700
rect 19230 17660 19270 17700
rect 19310 17660 19350 17700
rect 19390 17660 19430 17700
rect 19470 17660 19510 17700
rect 19550 17660 19590 17700
rect 19630 17660 19670 17700
rect 19710 17660 19750 17700
rect 19790 17660 19830 17700
rect 19870 17660 19910 17700
rect 19950 17660 19990 17700
rect 20030 17660 20070 17700
rect 20110 17660 20150 17700
rect 20190 17660 20230 17700
rect 20270 17660 20310 17700
rect 20350 17660 20390 17700
rect 20430 17660 20470 17700
rect 20510 17660 20550 17700
rect 20590 17660 20620 17700
rect 7280 17600 20620 17660
rect 7280 16790 19560 17600
rect 20370 16790 20620 17600
rect 7280 16740 20620 16790
rect 9620 16410 21160 16470
rect 9620 15720 10920 16410
rect 11750 15720 11950 16410
rect 12780 15720 12980 16410
rect 13810 15720 14040 16410
rect 14870 15720 15070 16410
rect 15900 15720 16100 16410
rect 16930 15720 17160 16410
rect 17990 15720 18190 16410
rect 19020 15720 19220 16410
rect 20050 15720 20280 16410
rect 21110 15720 21160 16410
rect 9620 15660 21160 15720
rect 9620 15620 9710 15660
rect 9750 15620 9790 15660
rect 9830 15620 9870 15660
rect 9910 15620 9950 15660
rect 9990 15620 10030 15660
rect 10070 15620 10110 15660
rect 10150 15620 10190 15660
rect 10230 15620 10270 15660
rect 10310 15620 10350 15660
rect 10390 15620 10430 15660
rect 10470 15620 10510 15660
rect 10550 15620 10590 15660
rect 10630 15620 10670 15660
rect 10710 15620 10750 15660
rect 10790 15620 10830 15660
rect 10870 15620 10910 15660
rect 10950 15620 10990 15660
rect 11030 15620 11070 15660
rect 11110 15620 11150 15660
rect 11190 15620 11230 15660
rect 11270 15620 11310 15660
rect 11350 15620 11390 15660
rect 11430 15620 11470 15660
rect 11510 15620 11550 15660
rect 11590 15620 11630 15660
rect 11670 15620 11710 15660
rect 11750 15620 11790 15660
rect 11830 15620 11870 15660
rect 11910 15620 11950 15660
rect 11990 15620 12030 15660
rect 12070 15620 12110 15660
rect 12150 15620 12190 15660
rect 12230 15620 12270 15660
rect 12310 15620 12350 15660
rect 12390 15620 12430 15660
rect 12470 15620 12510 15660
rect 12550 15620 12590 15660
rect 12630 15620 12670 15660
rect 12710 15620 12750 15660
rect 12790 15620 12830 15660
rect 12870 15620 12910 15660
rect 12950 15620 12990 15660
rect 13030 15620 13070 15660
rect 13110 15620 13150 15660
rect 13190 15620 13230 15660
rect 13270 15620 13310 15660
rect 13350 15620 13390 15660
rect 13430 15620 13470 15660
rect 13510 15620 13550 15660
rect 13590 15620 13630 15660
rect 13670 15620 13710 15660
rect 13750 15620 13790 15660
rect 13830 15620 13870 15660
rect 13910 15620 13950 15660
rect 13990 15620 14030 15660
rect 14070 15620 14110 15660
rect 14150 15620 14190 15660
rect 14230 15620 14270 15660
rect 14310 15620 14350 15660
rect 14390 15620 14430 15660
rect 14470 15620 14510 15660
rect 14550 15620 14590 15660
rect 14630 15620 14670 15660
rect 14710 15620 14750 15660
rect 14790 15620 14830 15660
rect 14870 15620 14910 15660
rect 14950 15620 14990 15660
rect 15030 15620 15070 15660
rect 15110 15620 15150 15660
rect 15190 15620 15230 15660
rect 15270 15620 15310 15660
rect 15350 15620 15390 15660
rect 15430 15620 15470 15660
rect 15510 15620 15550 15660
rect 15590 15620 15630 15660
rect 15670 15620 15710 15660
rect 15750 15620 15790 15660
rect 15830 15620 15870 15660
rect 15910 15620 15950 15660
rect 15990 15620 16030 15660
rect 16070 15620 16110 15660
rect 16150 15620 16190 15660
rect 16230 15620 16270 15660
rect 16310 15620 16350 15660
rect 16390 15620 16430 15660
rect 16470 15620 16510 15660
rect 16550 15620 16590 15660
rect 16630 15620 16670 15660
rect 16710 15620 16750 15660
rect 16790 15620 16830 15660
rect 16870 15620 16910 15660
rect 16950 15620 16990 15660
rect 17030 15620 17070 15660
rect 17110 15620 17150 15660
rect 17190 15620 17230 15660
rect 17270 15620 17310 15660
rect 17350 15620 17390 15660
rect 17430 15620 17470 15660
rect 17510 15620 17550 15660
rect 17590 15620 17630 15660
rect 17670 15620 17710 15660
rect 17750 15620 17790 15660
rect 17830 15620 17870 15660
rect 17910 15620 17950 15660
rect 17990 15620 18030 15660
rect 18070 15620 18110 15660
rect 18150 15620 18190 15660
rect 18230 15620 18270 15660
rect 18310 15620 18350 15660
rect 18390 15620 18430 15660
rect 18470 15620 18510 15660
rect 18550 15620 18590 15660
rect 18630 15620 18670 15660
rect 18710 15620 18750 15660
rect 18790 15620 18830 15660
rect 18870 15620 18910 15660
rect 18950 15620 18990 15660
rect 19030 15620 19070 15660
rect 19110 15620 19150 15660
rect 19190 15620 19230 15660
rect 19270 15620 19310 15660
rect 19350 15620 19390 15660
rect 19430 15620 19470 15660
rect 19510 15620 19550 15660
rect 19590 15620 19630 15660
rect 19670 15620 19710 15660
rect 19750 15620 19800 15660
rect 19840 15620 19880 15660
rect 19920 15620 19960 15660
rect 20000 15620 20040 15660
rect 20080 15620 20120 15660
rect 20160 15620 20200 15660
rect 20240 15620 20280 15660
rect 20320 15620 20370 15660
rect 20410 15620 20450 15660
rect 20490 15620 20530 15660
rect 20570 15620 20610 15660
rect 20650 15620 20690 15660
rect 20730 15620 20770 15660
rect 20810 15620 20850 15660
rect 20890 15620 20930 15660
rect 20970 15620 21010 15660
rect 21050 15620 21090 15660
rect 21130 15620 21160 15660
rect 9620 15610 21160 15620
rect 7420 15290 7510 15310
rect 7420 15230 7430 15290
rect 7500 15230 11260 15290
rect 7420 15210 7510 15230
rect 6740 15110 9830 15120
rect 6740 15050 9750 15110
rect 9810 15050 9830 15110
rect 6740 15040 9830 15050
rect 10060 15110 10630 15130
rect 10060 15080 10580 15110
rect 10060 15010 10100 15080
rect 10570 15070 10580 15080
rect 10620 15070 10630 15110
rect 10570 15050 10630 15070
rect 11200 15120 11260 15230
rect 11560 15120 11620 15130
rect 11200 15110 11620 15120
rect 12560 15110 12620 15130
rect 11200 15070 11570 15110
rect 11610 15070 11620 15110
rect 11200 15060 11620 15070
rect 11560 15050 11620 15060
rect 12510 15070 12570 15110
rect 12610 15070 12620 15110
rect 12510 15050 12620 15070
rect 10260 15020 10370 15030
rect 9940 15000 10120 15010
rect 9940 14960 10060 15000
rect 10100 14960 10120 15000
rect 9940 14950 10120 14960
rect 10260 14960 10280 15020
rect 10350 14960 10370 15020
rect 11300 15010 11360 15030
rect 12300 15010 12360 15030
rect 10260 14950 10370 14960
rect 10670 15000 10970 15010
rect 10670 14960 10820 15000
rect 10860 14960 10900 15000
rect 10940 14960 10970 15000
rect 10670 14950 10970 14960
rect 11080 15000 11310 15010
rect 11080 14960 11200 15000
rect 11240 14970 11310 15000
rect 11350 14970 11360 15010
rect 11240 14960 11360 14970
rect 11080 14950 11360 14960
rect 11660 15000 11960 15010
rect 11660 14960 11810 15000
rect 11850 14960 11890 15000
rect 11930 14960 11960 15000
rect 11660 14950 11960 14960
rect 12070 15000 12310 15010
rect 12070 14960 12190 15000
rect 12230 14970 12310 15000
rect 12350 14970 12360 15010
rect 12230 14960 12360 14970
rect 12070 14950 12360 14960
rect 10160 14350 10200 14360
rect 12510 14350 12560 15050
rect 13070 15010 13310 15030
rect 12660 15000 12960 15010
rect 12660 14960 12810 15000
rect 12850 14960 12890 15000
rect 12930 14960 12960 15000
rect 12660 14950 12960 14960
rect 13070 14970 13180 15010
rect 13220 14970 13260 15010
rect 13300 14970 13310 15010
rect 13070 14950 13310 14970
rect 13350 15010 13540 15030
rect 13350 14970 13360 15010
rect 13400 14970 13490 15010
rect 13530 14970 13540 15010
rect 13350 14950 13540 14970
rect 13690 15010 13880 15030
rect 13690 14970 13700 15010
rect 13740 14970 13830 15010
rect 13870 14970 13880 15010
rect 13690 14950 13880 14970
rect 14250 15010 14440 15030
rect 14250 14970 14260 15010
rect 14300 14970 14390 15010
rect 14430 14970 14440 15010
rect 14250 14950 14440 14970
rect 15250 15010 15500 15030
rect 15250 14970 15260 15010
rect 15300 14970 15450 15010
rect 15490 14970 15500 15010
rect 15250 14950 15500 14970
rect 17190 15020 17320 15030
rect 17190 14970 17250 15020
rect 17300 15010 17320 15020
rect 17380 15010 17450 15030
rect 17300 14970 17400 15010
rect 17440 14970 17450 15010
rect 17190 14960 17320 14970
rect 17380 14950 17450 14970
rect 20900 15020 22470 15030
rect 20900 14970 20960 15020
rect 21010 14970 22470 15020
rect 20900 14960 22470 14970
rect 9670 14340 21160 14350
rect 9670 14300 9700 14340
rect 9740 14300 9790 14340
rect 9830 14300 9870 14340
rect 9910 14300 9950 14340
rect 9990 14300 10030 14340
rect 10070 14300 10110 14340
rect 10150 14300 10190 14340
rect 10230 14300 10270 14340
rect 10310 14300 10350 14340
rect 10390 14300 10430 14340
rect 10470 14300 10510 14340
rect 10550 14300 10590 14340
rect 10630 14300 10670 14340
rect 10710 14300 10750 14340
rect 10790 14300 10830 14340
rect 10870 14300 10910 14340
rect 10950 14300 10990 14340
rect 11030 14300 11070 14340
rect 11110 14300 11150 14340
rect 11190 14300 11230 14340
rect 11270 14300 11310 14340
rect 11350 14300 11390 14340
rect 11430 14300 11470 14340
rect 11510 14300 11550 14340
rect 11590 14300 11630 14340
rect 11670 14300 11710 14340
rect 11750 14300 11790 14340
rect 11830 14300 11870 14340
rect 11910 14300 11950 14340
rect 11990 14300 12030 14340
rect 12070 14300 12110 14340
rect 12150 14300 12190 14340
rect 12230 14300 12270 14340
rect 12310 14300 12350 14340
rect 12390 14300 12430 14340
rect 12470 14300 12510 14340
rect 12550 14300 12590 14340
rect 12630 14300 12670 14340
rect 12710 14300 12750 14340
rect 12790 14300 12830 14340
rect 12870 14300 12910 14340
rect 12950 14300 12990 14340
rect 13030 14300 13070 14340
rect 13110 14300 13150 14340
rect 13230 14300 13270 14340
rect 13310 14300 13350 14340
rect 13390 14300 13430 14340
rect 13470 14300 13510 14340
rect 13550 14300 13590 14340
rect 13630 14300 13670 14340
rect 13710 14300 13750 14340
rect 13790 14300 13830 14340
rect 13870 14300 13910 14340
rect 13950 14300 13990 14340
rect 14030 14300 14070 14340
rect 14110 14300 14150 14340
rect 14190 14300 14230 14340
rect 14270 14300 14310 14340
rect 14350 14300 14390 14340
rect 14430 14300 14470 14340
rect 14510 14300 14550 14340
rect 14590 14300 14630 14340
rect 14670 14300 14710 14340
rect 14750 14300 14790 14340
rect 14830 14300 14870 14340
rect 14910 14300 14950 14340
rect 14990 14300 15030 14340
rect 15070 14300 15110 14340
rect 15150 14300 15190 14340
rect 15230 14300 15270 14340
rect 15310 14300 15350 14340
rect 15390 14300 15430 14340
rect 15470 14300 15510 14340
rect 15550 14300 15590 14340
rect 15630 14300 15670 14340
rect 15710 14300 15750 14340
rect 15790 14300 15830 14340
rect 15870 14300 15910 14340
rect 15950 14300 15990 14340
rect 16030 14300 16070 14340
rect 16110 14300 16150 14340
rect 16190 14300 16230 14340
rect 16270 14300 16310 14340
rect 16350 14300 16390 14340
rect 16430 14300 16470 14340
rect 16510 14300 16550 14340
rect 16590 14300 16630 14340
rect 16670 14300 16710 14340
rect 16750 14300 16790 14340
rect 16830 14300 16870 14340
rect 16910 14300 16950 14340
rect 16990 14300 17030 14340
rect 17070 14300 17110 14340
rect 17150 14300 17190 14340
rect 17230 14300 17270 14340
rect 17310 14300 17350 14340
rect 17390 14300 17430 14340
rect 17470 14300 17510 14340
rect 17550 14300 17590 14340
rect 17630 14300 17670 14340
rect 17710 14300 17750 14340
rect 17790 14300 17830 14340
rect 17870 14300 17910 14340
rect 17950 14300 17990 14340
rect 18030 14300 18070 14340
rect 18110 14300 18150 14340
rect 18190 14300 18230 14340
rect 18270 14300 18310 14340
rect 18350 14300 18390 14340
rect 18430 14300 18470 14340
rect 18510 14300 18550 14340
rect 18590 14300 18630 14340
rect 18670 14300 18710 14340
rect 18750 14300 18790 14340
rect 18830 14300 18870 14340
rect 18910 14300 18950 14340
rect 18990 14300 19030 14340
rect 19070 14300 19110 14340
rect 19150 14300 19190 14340
rect 19230 14300 19270 14340
rect 19310 14300 19350 14340
rect 19390 14300 19430 14340
rect 19470 14300 19510 14340
rect 19550 14300 19590 14340
rect 19630 14300 19670 14340
rect 19710 14300 19750 14340
rect 19790 14300 19830 14340
rect 19870 14300 19910 14340
rect 19950 14300 19990 14340
rect 20030 14300 20070 14340
rect 20110 14300 20150 14340
rect 20190 14300 20230 14340
rect 20270 14300 20310 14340
rect 20350 14300 20390 14340
rect 20430 14300 20470 14340
rect 20510 14300 20550 14340
rect 20590 14300 20630 14340
rect 20670 14300 20710 14340
rect 20750 14300 20790 14340
rect 20830 14300 20870 14340
rect 20910 14300 20950 14340
rect 20990 14300 21030 14340
rect 21070 14300 21160 14340
rect 9670 14290 21160 14300
rect 7280 14260 21160 14290
rect 7280 14200 8430 14260
rect 8500 14240 21160 14260
rect 8500 14200 9910 14240
rect 7280 13430 9910 14200
rect 10720 13430 10940 14240
rect 11750 13430 11970 14240
rect 12780 13430 12980 14240
rect 13790 13430 21160 14240
rect 7280 13370 21160 13430
rect 7280 13330 7320 13370
rect 7360 13330 7400 13370
rect 7440 13330 7480 13370
rect 7520 13330 7560 13370
rect 7600 13330 7640 13370
rect 7680 13330 7720 13370
rect 7760 13330 7800 13370
rect 7840 13330 7880 13370
rect 7920 13330 7960 13370
rect 8000 13330 8040 13370
rect 8080 13330 8120 13370
rect 8160 13330 8200 13370
rect 8240 13330 8280 13370
rect 8320 13330 8360 13370
rect 8400 13330 8440 13370
rect 8480 13330 8520 13370
rect 8560 13330 8600 13370
rect 8640 13330 8680 13370
rect 8720 13330 8760 13370
rect 8800 13330 8840 13370
rect 8880 13330 8920 13370
rect 8960 13330 9000 13370
rect 9040 13330 9080 13370
rect 9120 13330 9160 13370
rect 9200 13330 9240 13370
rect 9280 13330 9320 13370
rect 9360 13330 9400 13370
rect 9440 13330 9480 13370
rect 9520 13330 9560 13370
rect 9600 13330 9640 13370
rect 9680 13330 9720 13370
rect 9760 13330 9800 13370
rect 9840 13330 9890 13370
rect 9930 13330 9970 13370
rect 10010 13330 10050 13370
rect 10090 13330 10130 13370
rect 10170 13330 10210 13370
rect 10250 13330 10290 13370
rect 10330 13330 10370 13370
rect 10410 13330 10450 13370
rect 10490 13330 10530 13370
rect 10570 13330 10610 13370
rect 10650 13330 10690 13370
rect 10730 13330 10770 13370
rect 10810 13330 10850 13370
rect 10890 13330 10930 13370
rect 10970 13330 11010 13370
rect 11050 13330 11090 13370
rect 11130 13330 11170 13370
rect 11210 13330 11250 13370
rect 11290 13330 11330 13370
rect 11370 13330 11410 13370
rect 11450 13330 11490 13370
rect 11530 13330 11570 13370
rect 11610 13330 11650 13370
rect 11690 13330 11730 13370
rect 11770 13330 11810 13370
rect 11850 13330 11890 13370
rect 11930 13330 11970 13370
rect 12010 13330 12050 13370
rect 12090 13330 12130 13370
rect 12170 13330 12210 13370
rect 12250 13330 12290 13370
rect 12330 13330 12370 13370
rect 12410 13330 12450 13370
rect 12490 13330 12530 13370
rect 12570 13330 12610 13370
rect 12650 13330 12690 13370
rect 12730 13330 12770 13370
rect 12810 13330 12850 13370
rect 12890 13330 12930 13370
rect 12970 13330 13010 13370
rect 13050 13330 13090 13370
rect 13130 13330 13170 13370
rect 13210 13330 13250 13370
rect 13290 13330 13330 13370
rect 13400 13330 13440 13370
rect 13480 13330 13520 13370
rect 13560 13330 13600 13370
rect 13640 13330 13680 13370
rect 13720 13330 13760 13370
rect 13800 13330 13840 13370
rect 13880 13330 13920 13370
rect 13960 13330 14000 13370
rect 14040 13330 14080 13370
rect 14120 13330 14160 13370
rect 14200 13330 14240 13370
rect 14280 13330 14320 13370
rect 14360 13330 14400 13370
rect 14440 13330 14480 13370
rect 14520 13330 14560 13370
rect 14600 13330 14640 13370
rect 14680 13330 14720 13370
rect 14760 13330 14800 13370
rect 14840 13330 14880 13370
rect 14920 13330 14960 13370
rect 15000 13330 15040 13370
rect 15080 13330 15120 13370
rect 15160 13330 15200 13370
rect 15240 13330 15280 13370
rect 15320 13330 15360 13370
rect 15400 13330 15440 13370
rect 15480 13330 15520 13370
rect 15560 13330 15600 13370
rect 15640 13330 15680 13370
rect 15720 13330 15760 13370
rect 15800 13330 15840 13370
rect 15880 13330 15920 13370
rect 15960 13330 16000 13370
rect 16040 13330 16080 13370
rect 16120 13330 16160 13370
rect 16200 13330 16240 13370
rect 16280 13330 16320 13370
rect 16360 13330 16400 13370
rect 16440 13330 16480 13370
rect 16520 13330 16560 13370
rect 16600 13330 16640 13370
rect 16680 13330 16720 13370
rect 16760 13330 16800 13370
rect 16840 13330 16880 13370
rect 16920 13330 16960 13370
rect 17000 13330 17040 13370
rect 17080 13330 17120 13370
rect 17160 13330 17200 13370
rect 17240 13330 17280 13370
rect 17320 13330 17360 13370
rect 17400 13330 17440 13370
rect 17480 13330 17520 13370
rect 17560 13330 17600 13370
rect 17640 13330 17680 13370
rect 17720 13330 17760 13370
rect 17800 13330 17840 13370
rect 17880 13330 17920 13370
rect 17960 13330 18000 13370
rect 18040 13330 18080 13370
rect 18120 13330 18160 13370
rect 18200 13330 18240 13370
rect 18280 13330 18320 13370
rect 18360 13330 18400 13370
rect 18440 13330 18480 13370
rect 18520 13330 18560 13370
rect 18600 13330 18640 13370
rect 18680 13330 18720 13370
rect 18760 13330 18800 13370
rect 18840 13330 18880 13370
rect 18920 13330 18960 13370
rect 19000 13330 19040 13370
rect 19080 13330 19120 13370
rect 19160 13330 19200 13370
rect 19240 13330 19280 13370
rect 19320 13330 19360 13370
rect 19400 13330 19440 13370
rect 19480 13330 19520 13370
rect 19560 13330 19600 13370
rect 19640 13330 19680 13370
rect 19720 13330 19760 13370
rect 19800 13330 19840 13370
rect 19880 13330 19920 13370
rect 19960 13330 20000 13370
rect 20040 13330 20080 13370
rect 20120 13330 20160 13370
rect 20200 13330 20240 13370
rect 20280 13330 20320 13370
rect 20360 13330 20400 13370
rect 20440 13330 20480 13370
rect 20520 13330 20560 13370
rect 20600 13330 20640 13370
rect 20680 13330 20720 13370
rect 20760 13330 20800 13370
rect 20840 13330 20880 13370
rect 20920 13330 20960 13370
rect 21000 13330 21040 13370
rect 21080 13330 21160 13370
rect 7280 13320 21160 13330
rect 5610 12720 5730 12730
rect 5610 12710 7350 12720
rect 5610 12650 7270 12710
rect 7330 12650 7350 12710
rect 5610 12640 7350 12650
rect 7460 12710 7870 12720
rect 7460 12700 7700 12710
rect 7460 12660 7570 12700
rect 7610 12660 7700 12700
rect 7460 12650 7700 12660
rect 7760 12700 7870 12710
rect 7760 12660 7820 12700
rect 7860 12660 7870 12700
rect 8170 12710 8380 12720
rect 8170 12670 8320 12710
rect 8360 12670 8380 12710
rect 8170 12660 8380 12670
rect 7760 12650 7870 12660
rect 7460 12640 7870 12650
rect 7570 12600 7670 12610
rect 8070 12600 8130 12620
rect 7570 12540 7590 12600
rect 7650 12560 8080 12600
rect 8120 12560 8130 12600
rect 7650 12540 8130 12560
rect 8320 12590 8380 12660
rect 8440 12710 8490 13320
rect 9660 13150 9810 13170
rect 9660 13090 9670 13150
rect 9740 13090 9810 13150
rect 9660 13070 9810 13090
rect 9760 12720 9810 13070
rect 8440 12690 8620 12710
rect 8440 12650 8570 12690
rect 8610 12650 8620 12690
rect 8440 12630 8620 12650
rect 8800 12700 9000 12720
rect 8800 12660 8870 12700
rect 8910 12660 8950 12700
rect 8990 12660 9000 12700
rect 8800 12640 9000 12660
rect 9040 12700 9260 12720
rect 9040 12660 9070 12700
rect 9110 12660 9210 12700
rect 9250 12660 9260 12700
rect 9040 12640 9260 12660
rect 9300 12700 9510 12720
rect 9300 12660 9330 12700
rect 9370 12660 9460 12700
rect 9500 12660 9510 12700
rect 9300 12640 9510 12660
rect 9550 12700 9680 12720
rect 9550 12660 9580 12700
rect 9620 12660 9680 12700
rect 9550 12640 9680 12660
rect 8700 12590 8770 12600
rect 8320 12580 8770 12590
rect 8320 12540 8720 12580
rect 8760 12540 8770 12580
rect 7570 12530 7670 12540
rect 8320 12530 8770 12540
rect 8700 12520 8770 12530
rect 9640 12390 9680 12640
rect 9760 12710 9930 12720
rect 9760 12670 9860 12710
rect 9900 12670 9930 12710
rect 9760 12660 9930 12670
rect 10040 12710 10220 12720
rect 10040 12670 10160 12710
rect 10200 12670 10220 12710
rect 10040 12660 10220 12670
rect 10260 12700 10300 13320
rect 10410 12700 10470 12720
rect 10260 12660 10420 12700
rect 10460 12660 10470 12700
rect 10770 12710 11070 12720
rect 10770 12670 10920 12710
rect 10960 12670 11000 12710
rect 11040 12670 11070 12710
rect 10770 12660 11070 12670
rect 11180 12710 11460 12720
rect 11180 12670 11300 12710
rect 11340 12700 11460 12710
rect 11340 12670 11410 12700
rect 11180 12660 11410 12670
rect 11450 12660 11460 12700
rect 11760 12710 12060 12720
rect 11760 12670 11910 12710
rect 11950 12670 11990 12710
rect 12030 12670 12060 12710
rect 11760 12660 12060 12670
rect 12170 12710 12460 12720
rect 12170 12670 12290 12710
rect 12330 12700 12460 12710
rect 12330 12670 12410 12700
rect 12170 12660 12410 12670
rect 12450 12660 12460 12700
rect 12760 12710 13060 12720
rect 12760 12670 12910 12710
rect 12950 12670 12990 12710
rect 13030 12670 13060 12710
rect 12760 12660 13060 12670
rect 13170 12700 13410 12720
rect 13170 12660 13280 12700
rect 13320 12660 13360 12700
rect 13400 12660 13410 12700
rect 9760 12550 9810 12660
rect 10160 12600 10200 12660
rect 10410 12640 10470 12660
rect 11400 12640 11460 12660
rect 12400 12640 12460 12660
rect 13170 12640 13410 12660
rect 13450 12700 13640 12720
rect 13450 12660 13460 12700
rect 13500 12660 13590 12700
rect 13630 12660 13640 12700
rect 13450 12640 13640 12660
rect 13790 12700 13980 12720
rect 13790 12660 13800 12700
rect 13840 12660 13930 12700
rect 13970 12660 13980 12700
rect 13790 12640 13980 12660
rect 14350 12700 14540 12720
rect 14350 12660 14360 12700
rect 14400 12660 14490 12700
rect 14530 12660 14540 12700
rect 14350 12640 14540 12660
rect 15350 12700 15600 12720
rect 15350 12660 15360 12700
rect 15400 12660 15550 12700
rect 15590 12660 15600 12700
rect 15350 12640 15600 12660
rect 17290 12700 17420 12710
rect 17480 12700 17550 12720
rect 17290 12650 17350 12700
rect 17400 12660 17500 12700
rect 17540 12660 17550 12700
rect 17400 12650 17420 12660
rect 17290 12640 17420 12650
rect 17480 12640 17550 12660
rect 21000 12700 22040 12710
rect 21000 12650 21060 12700
rect 21110 12650 22040 12700
rect 21000 12640 22040 12650
rect 10670 12600 10730 12620
rect 10160 12560 10680 12600
rect 10720 12560 10730 12600
rect 9740 12530 9830 12550
rect 10670 12540 10730 12560
rect 11270 12610 11360 12630
rect 11660 12610 11720 12620
rect 11270 12550 11280 12610
rect 11350 12600 11720 12610
rect 11350 12560 11670 12600
rect 11710 12560 11720 12600
rect 11350 12550 11720 12560
rect 11270 12530 11360 12550
rect 11660 12540 11720 12550
rect 12660 12600 12720 12620
rect 12660 12560 12670 12600
rect 12710 12560 12720 12600
rect 12660 12540 12720 12560
rect 9740 12470 9750 12530
rect 9820 12470 9830 12530
rect 9740 12450 9830 12470
rect 12660 12390 12710 12540
rect 9640 12350 12710 12390
rect 9730 12050 21160 12060
rect 9730 12010 9810 12050
rect 9850 12010 9890 12050
rect 9930 12010 9970 12050
rect 10010 12010 10050 12050
rect 10090 12010 10130 12050
rect 10170 12010 10210 12050
rect 10250 12010 10290 12050
rect 10330 12010 10370 12050
rect 10410 12010 10450 12050
rect 10490 12010 10530 12050
rect 10570 12010 10610 12050
rect 10650 12010 10690 12050
rect 10730 12010 10770 12050
rect 10810 12010 10850 12050
rect 10890 12010 10930 12050
rect 10970 12010 11010 12050
rect 11050 12010 11090 12050
rect 11130 12010 11170 12050
rect 11210 12010 11250 12050
rect 11290 12010 11330 12050
rect 11370 12010 11410 12050
rect 11450 12010 11490 12050
rect 11530 12010 11570 12050
rect 11610 12010 11650 12050
rect 11690 12010 11730 12050
rect 11770 12010 11810 12050
rect 11850 12010 11890 12050
rect 11930 12010 11970 12050
rect 12010 12010 12050 12050
rect 12090 12010 12130 12050
rect 12170 12010 12210 12050
rect 12250 12010 12290 12050
rect 12330 12010 12370 12050
rect 12410 12010 12450 12050
rect 12490 12010 12530 12050
rect 12570 12010 12610 12050
rect 12650 12010 12690 12050
rect 12730 12010 12770 12050
rect 12810 12010 12850 12050
rect 12890 12010 12930 12050
rect 12970 12010 13010 12050
rect 13050 12010 13090 12050
rect 13130 12010 13170 12050
rect 13210 12010 13250 12050
rect 13290 12010 13330 12050
rect 13440 12010 13480 12050
rect 13520 12010 13560 12050
rect 13600 12010 13640 12050
rect 13680 12010 13720 12050
rect 13760 12010 13800 12050
rect 13840 12010 13880 12050
rect 13920 12010 13960 12050
rect 14000 12010 14040 12050
rect 14080 12010 14120 12050
rect 14160 12010 14200 12050
rect 14240 12010 14280 12050
rect 14320 12010 14360 12050
rect 14400 12010 14440 12050
rect 14480 12010 14520 12050
rect 14560 12010 14600 12050
rect 14640 12010 14680 12050
rect 14720 12010 14760 12050
rect 14800 12010 14840 12050
rect 14880 12010 14920 12050
rect 14960 12010 15000 12050
rect 15040 12010 15080 12050
rect 15120 12010 15160 12050
rect 15200 12010 15240 12050
rect 15280 12010 15320 12050
rect 15360 12010 15400 12050
rect 15440 12010 15480 12050
rect 15520 12010 15560 12050
rect 15600 12010 15640 12050
rect 15680 12010 15720 12050
rect 15760 12010 15800 12050
rect 15840 12010 15880 12050
rect 15920 12010 15960 12050
rect 16000 12010 16040 12050
rect 16080 12010 16120 12050
rect 16160 12010 16200 12050
rect 16240 12010 16280 12050
rect 16320 12010 16360 12050
rect 16400 12010 16440 12050
rect 16480 12010 16520 12050
rect 16560 12010 16600 12050
rect 16640 12010 16680 12050
rect 16720 12010 16760 12050
rect 16800 12010 16840 12050
rect 16880 12010 16920 12050
rect 16960 12010 17000 12050
rect 17040 12010 17080 12050
rect 17120 12010 17160 12050
rect 17200 12010 17240 12050
rect 17280 12010 17320 12050
rect 17360 12010 17400 12050
rect 17440 12010 17480 12050
rect 17520 12010 17560 12050
rect 17600 12010 17640 12050
rect 17680 12010 17720 12050
rect 17760 12010 17800 12050
rect 17840 12010 17880 12050
rect 17920 12010 17960 12050
rect 18000 12010 18040 12050
rect 18080 12010 18120 12050
rect 18160 12010 18200 12050
rect 18240 12010 18280 12050
rect 18320 12010 18360 12050
rect 18400 12010 18440 12050
rect 18480 12010 18520 12050
rect 18560 12010 18600 12050
rect 18640 12010 18680 12050
rect 18720 12010 18760 12050
rect 18800 12010 18840 12050
rect 18880 12010 18920 12050
rect 18960 12010 19000 12050
rect 19040 12010 19080 12050
rect 19120 12010 19160 12050
rect 19200 12010 19240 12050
rect 19280 12010 19320 12050
rect 19360 12010 19400 12050
rect 19440 12010 19480 12050
rect 19520 12010 19560 12050
rect 19600 12010 19640 12050
rect 19680 12010 19720 12050
rect 19760 12010 19800 12050
rect 19840 12010 19890 12050
rect 19930 12010 19970 12050
rect 20010 12010 20050 12050
rect 20090 12010 20130 12050
rect 20170 12010 20210 12050
rect 20250 12010 20290 12050
rect 20330 12010 20370 12050
rect 20410 12010 20460 12050
rect 20500 12010 20540 12050
rect 20580 12010 20620 12050
rect 20660 12010 20700 12050
rect 20740 12010 20780 12050
rect 20820 12010 20860 12050
rect 20900 12010 20940 12050
rect 20980 12010 21020 12050
rect 21060 12010 21160 12050
rect 7280 12000 21160 12010
rect 7280 11960 7330 12000
rect 7370 11960 7410 12000
rect 7450 11960 7490 12000
rect 7530 11960 7570 12000
rect 7610 11960 7650 12000
rect 7690 11960 7730 12000
rect 7770 11960 7810 12000
rect 7850 11960 7890 12000
rect 7930 11960 7970 12000
rect 8010 11960 8050 12000
rect 8090 11960 8130 12000
rect 8170 11960 8210 12000
rect 8250 11960 8290 12000
rect 8330 11960 8370 12000
rect 8410 11960 8450 12000
rect 8490 11960 8530 12000
rect 8570 11960 8610 12000
rect 8650 11960 8690 12000
rect 8730 11960 8770 12000
rect 8810 11960 8850 12000
rect 8890 11960 8930 12000
rect 8970 11960 9010 12000
rect 9050 11960 9090 12000
rect 9130 11960 9170 12000
rect 9210 11960 9250 12000
rect 9290 11960 9330 12000
rect 9370 11960 9410 12000
rect 9450 11960 9490 12000
rect 9530 11960 9570 12000
rect 9610 11960 9650 12000
rect 9690 11960 9730 12000
rect 9770 11960 21160 12000
rect 7280 11860 21160 11960
rect 7280 11410 14040 11860
rect 7280 11370 7720 11410
rect 7760 11370 7800 11410
rect 7840 11370 7880 11410
rect 7920 11370 7960 11410
rect 8000 11370 8040 11410
rect 8080 11370 8120 11410
rect 8160 11370 8200 11410
rect 8240 11370 8280 11410
rect 8320 11370 8360 11410
rect 8400 11370 8440 11410
rect 8480 11370 8520 11410
rect 8560 11370 14040 11410
rect 7280 11360 14040 11370
rect 7280 11330 7720 11360
rect 7280 11290 7670 11330
rect 7710 11290 7720 11330
rect 7280 11250 7720 11290
rect 7280 11210 7670 11250
rect 7710 11210 7720 11250
rect 7280 11170 7720 11210
rect 7280 11130 7670 11170
rect 7710 11130 7720 11170
rect 7280 11090 7720 11130
rect 7280 11050 7330 11090
rect 7370 11050 7410 11090
rect 7450 11050 7490 11090
rect 7530 11050 7570 11090
rect 7610 11050 7650 11090
rect 7690 11050 7720 11090
rect 7280 11040 7720 11050
rect 8540 11330 14040 11360
rect 8540 11290 8550 11330
rect 8590 11290 14040 11330
rect 8540 11250 14040 11290
rect 8540 11210 8550 11250
rect 8590 11210 14040 11250
rect 8540 11170 14040 11210
rect 14870 11170 15070 11860
rect 15900 11170 16100 11860
rect 16930 11170 17160 11860
rect 17990 11170 18190 11860
rect 19020 11170 19220 11860
rect 20050 11170 20280 11860
rect 21110 11170 21160 11860
rect 8540 11130 8550 11170
rect 8590 11130 21160 11170
rect 8540 11090 21160 11130
rect 8540 11050 8610 11090
rect 8650 11050 8690 11090
rect 8730 11050 8770 11090
rect 8810 11050 8850 11090
rect 8890 11050 8930 11090
rect 8970 11050 9010 11090
rect 9050 11050 9090 11090
rect 9130 11050 9170 11090
rect 9210 11050 9250 11090
rect 9290 11050 9330 11090
rect 9370 11050 9410 11090
rect 9450 11050 9490 11090
rect 9530 11050 9570 11090
rect 9610 11050 9650 11090
rect 9690 11050 9730 11090
rect 9770 11050 21160 11090
rect 8540 11040 21160 11050
rect 9730 11000 9810 11040
rect 9850 11000 9890 11040
rect 9930 11000 9970 11040
rect 10010 11000 10050 11040
rect 10090 11000 10130 11040
rect 10170 11000 10210 11040
rect 10250 11000 10290 11040
rect 10330 11000 10370 11040
rect 10410 11000 10450 11040
rect 10490 11000 10530 11040
rect 10570 11000 10610 11040
rect 10650 11000 10690 11040
rect 10730 11000 10770 11040
rect 10810 11000 10850 11040
rect 10890 11000 10930 11040
rect 10970 11000 11010 11040
rect 11050 11000 11090 11040
rect 11130 11000 11170 11040
rect 11210 11000 11250 11040
rect 11290 11000 11330 11040
rect 11370 11000 11410 11040
rect 11450 11000 11490 11040
rect 11530 11000 11570 11040
rect 11610 11000 11650 11040
rect 11690 11000 11730 11040
rect 11770 11000 11810 11040
rect 11850 11000 11890 11040
rect 11930 11000 11970 11040
rect 12010 11000 12050 11040
rect 12090 11000 12130 11040
rect 12170 11000 12210 11040
rect 12250 11000 12290 11040
rect 12330 11000 12370 11040
rect 12410 11000 12450 11040
rect 12490 11000 12530 11040
rect 12570 11000 12610 11040
rect 12650 11000 12690 11040
rect 12730 11000 12770 11040
rect 12810 11000 12850 11040
rect 12890 11000 12930 11040
rect 12970 11000 13010 11040
rect 13050 11000 13090 11040
rect 13130 11000 13170 11040
rect 13210 11000 13250 11040
rect 13290 11000 13330 11040
rect 13410 11000 13450 11040
rect 13490 11000 13530 11040
rect 13570 11000 13610 11040
rect 13650 11000 13690 11040
rect 13730 11000 13770 11040
rect 13810 11000 13850 11040
rect 13890 11000 13930 11040
rect 13970 11000 14010 11040
rect 14050 11000 14090 11040
rect 14130 11000 14170 11040
rect 14210 11000 14250 11040
rect 14290 11000 14330 11040
rect 14370 11000 14410 11040
rect 14450 11000 14490 11040
rect 14530 11000 14570 11040
rect 14610 11000 14650 11040
rect 14690 11000 14730 11040
rect 14770 11000 14810 11040
rect 14850 11000 14890 11040
rect 14930 11000 14970 11040
rect 15010 11000 15050 11040
rect 15090 11000 15130 11040
rect 15170 11000 15210 11040
rect 15250 11000 15290 11040
rect 15330 11000 15370 11040
rect 15410 11000 15450 11040
rect 15490 11000 15530 11040
rect 15570 11000 15610 11040
rect 15650 11000 15690 11040
rect 15730 11000 15770 11040
rect 15810 11000 15850 11040
rect 15890 11000 15930 11040
rect 15970 11000 16010 11040
rect 16050 11000 16090 11040
rect 16130 11000 16170 11040
rect 16210 11000 16250 11040
rect 16290 11000 16330 11040
rect 16370 11000 16410 11040
rect 16450 11000 16490 11040
rect 16530 11000 16570 11040
rect 16610 11000 16650 11040
rect 16690 11000 16730 11040
rect 16770 11000 16810 11040
rect 16850 11000 16890 11040
rect 16930 11000 16970 11040
rect 17010 11000 17050 11040
rect 17090 11000 17130 11040
rect 17170 11000 17210 11040
rect 17250 11000 17290 11040
rect 17330 11000 17370 11040
rect 17410 11000 17450 11040
rect 17490 11000 17530 11040
rect 17570 11000 17610 11040
rect 17650 11000 17690 11040
rect 17730 11000 17770 11040
rect 17810 11000 17850 11040
rect 17890 11000 17930 11040
rect 17970 11000 18010 11040
rect 18050 11000 18090 11040
rect 18130 11000 18170 11040
rect 18210 11000 18250 11040
rect 18290 11000 18330 11040
rect 18370 11000 18410 11040
rect 18450 11000 18490 11040
rect 18530 11000 18570 11040
rect 18610 11000 18650 11040
rect 18690 11000 18730 11040
rect 18770 11000 18810 11040
rect 18850 11000 18890 11040
rect 18930 11000 18970 11040
rect 19010 11000 19050 11040
rect 19090 11000 19130 11040
rect 19170 11000 19210 11040
rect 19250 11000 19290 11040
rect 19330 11000 19370 11040
rect 19410 11000 19450 11040
rect 19490 11000 19540 11040
rect 19580 11000 19620 11040
rect 19660 11000 19700 11040
rect 19740 11000 19780 11040
rect 19820 11000 19860 11040
rect 19900 11000 19940 11040
rect 19980 11000 20020 11040
rect 20060 11000 20110 11040
rect 20150 11000 20190 11040
rect 20230 11000 20270 11040
rect 20310 11000 20350 11040
rect 20390 11000 20430 11040
rect 20470 11000 20510 11040
rect 20550 11000 20590 11040
rect 20630 11000 20670 11040
rect 20710 11000 20750 11040
rect 20790 11000 20830 11040
rect 20870 11000 20910 11040
rect 20950 11000 20990 11040
rect 21030 11000 21070 11040
rect 21110 11000 21160 11040
rect 9730 10990 21160 11000
rect 7590 10950 7690 10960
rect 7590 10890 7610 10950
rect 7670 10940 7690 10950
rect 8120 10940 8180 10960
rect 7670 10900 8130 10940
rect 8170 10900 8180 10940
rect 7670 10890 7690 10900
rect 7590 10880 7690 10890
rect 8120 10880 8180 10900
rect 8330 10940 8530 10950
rect 8330 10900 8350 10940
rect 8390 10900 8530 10940
rect 8330 10890 8530 10900
rect 5380 10410 7350 10420
rect 5380 10350 7270 10410
rect 7330 10350 7350 10410
rect 7600 10390 7670 10880
rect 7840 10850 7920 10870
rect 7840 10790 7850 10850
rect 7910 10790 7920 10850
rect 7840 10770 7920 10790
rect 8470 10530 8530 10890
rect 9630 10840 9740 10860
rect 9630 10780 9650 10840
rect 9720 10780 9830 10840
rect 9630 10760 9740 10780
rect 9770 10690 9830 10780
rect 9770 10680 9930 10690
rect 9770 10640 9860 10680
rect 9900 10640 9930 10680
rect 9770 10630 9930 10640
rect 8790 10530 8860 10540
rect 8470 10520 8860 10530
rect 8470 10480 8810 10520
rect 8850 10480 8860 10520
rect 11280 10530 11370 10550
rect 10670 10490 10730 10510
rect 8470 10470 8860 10480
rect 8790 10460 8860 10470
rect 10160 10450 10680 10490
rect 10720 10450 10730 10490
rect 11280 10470 11290 10530
rect 11360 10490 11370 10530
rect 11660 10490 11720 10510
rect 11360 10470 11670 10490
rect 11280 10450 11670 10470
rect 11710 10450 11720 10490
rect 5380 10340 7350 10350
rect 7460 10380 7670 10390
rect 7460 10340 7610 10380
rect 7650 10340 7670 10380
rect 7460 10330 7670 10340
rect 8540 10410 8710 10430
rect 8540 10370 8660 10410
rect 8700 10370 8710 10410
rect 8540 10350 8710 10370
rect 8890 10400 9090 10420
rect 8890 10360 8960 10400
rect 9000 10360 9040 10400
rect 9080 10360 9090 10400
rect 8540 9730 8590 10350
rect 8890 10340 9090 10360
rect 9130 10400 9350 10420
rect 9130 10360 9160 10400
rect 9200 10360 9300 10400
rect 9340 10360 9350 10400
rect 9130 10340 9350 10360
rect 9390 10400 9600 10420
rect 9390 10360 9420 10400
rect 9460 10360 9550 10400
rect 9590 10360 9600 10400
rect 9390 10340 9600 10360
rect 9640 10410 9720 10420
rect 9770 10410 9880 10430
rect 9640 10400 9790 10410
rect 9640 10360 9670 10400
rect 9710 10360 9790 10400
rect 9640 10350 9790 10360
rect 9860 10350 9880 10410
rect 10160 10390 10200 10450
rect 10670 10430 10730 10450
rect 11660 10430 11720 10450
rect 12280 10500 12370 10520
rect 12660 10500 12720 10510
rect 12280 10440 12290 10500
rect 12360 10490 12720 10500
rect 12360 10450 12670 10490
rect 12710 10450 12720 10490
rect 12360 10440 12720 10450
rect 12280 10420 12370 10440
rect 12660 10430 12720 10440
rect 10410 10390 10470 10410
rect 11400 10390 11460 10410
rect 12400 10390 12460 10410
rect 13170 10390 13400 10410
rect 9640 10340 9720 10350
rect 9770 10330 9880 10350
rect 10040 10380 10220 10390
rect 10040 10340 10160 10380
rect 10200 10340 10220 10380
rect 10040 10330 10220 10340
rect 10260 10350 10420 10390
rect 10460 10350 10470 10390
rect 10260 9730 10300 10350
rect 10410 10330 10470 10350
rect 10770 10380 11070 10390
rect 10770 10340 10920 10380
rect 10960 10340 11000 10380
rect 11040 10340 11070 10380
rect 10770 10330 11070 10340
rect 11180 10380 11410 10390
rect 11180 10340 11300 10380
rect 11340 10350 11410 10380
rect 11450 10350 11460 10390
rect 11340 10340 11460 10350
rect 11180 10330 11460 10340
rect 11760 10380 12060 10390
rect 11760 10340 11910 10380
rect 11950 10340 11990 10380
rect 12030 10340 12060 10380
rect 11760 10330 12060 10340
rect 12170 10380 12410 10390
rect 12170 10340 12290 10380
rect 12330 10350 12410 10380
rect 12450 10350 12460 10390
rect 12330 10340 12460 10350
rect 12170 10330 12460 10340
rect 12760 10380 13060 10390
rect 12760 10340 12910 10380
rect 12950 10340 12990 10380
rect 13030 10340 13060 10380
rect 12760 10330 13060 10340
rect 13170 10350 13270 10390
rect 13310 10350 13350 10390
rect 13390 10350 13400 10390
rect 13170 10330 13400 10350
rect 13440 10390 13630 10410
rect 13440 10350 13450 10390
rect 13490 10350 13580 10390
rect 13620 10350 13630 10390
rect 13440 10330 13630 10350
rect 13780 10390 13970 10410
rect 13780 10350 13790 10390
rect 13830 10350 13920 10390
rect 13960 10350 13970 10390
rect 13780 10330 13970 10350
rect 14340 10390 14530 10410
rect 14340 10350 14350 10390
rect 14390 10350 14480 10390
rect 14520 10350 14530 10390
rect 14340 10330 14530 10350
rect 15340 10390 15590 10410
rect 15340 10350 15350 10390
rect 15390 10350 15540 10390
rect 15580 10350 15590 10390
rect 15340 10330 15590 10350
rect 17280 10400 17410 10410
rect 17280 10350 17340 10400
rect 17390 10390 17410 10400
rect 17470 10390 17540 10410
rect 17390 10350 17490 10390
rect 17530 10350 17540 10390
rect 17280 10340 17410 10350
rect 17470 10330 17540 10350
rect 20990 10400 21640 10410
rect 20990 10350 21050 10400
rect 21100 10350 21640 10400
rect 20990 10340 21640 10350
rect 7280 9720 7790 9730
rect 7280 9680 7320 9720
rect 7360 9680 7400 9720
rect 7440 9680 7480 9720
rect 7520 9680 7560 9720
rect 7600 9680 7640 9720
rect 7680 9680 7720 9720
rect 7760 9680 7790 9720
rect 7280 9650 7790 9680
rect 8470 9720 21160 9730
rect 8470 9680 8520 9720
rect 8560 9680 8600 9720
rect 8640 9680 8680 9720
rect 8720 9680 8760 9720
rect 8800 9680 8840 9720
rect 8880 9680 8920 9720
rect 8960 9680 9000 9720
rect 9040 9680 9080 9720
rect 9120 9680 9160 9720
rect 9200 9680 9240 9720
rect 9280 9680 9320 9720
rect 9360 9680 9400 9720
rect 9440 9680 9480 9720
rect 9520 9680 9560 9720
rect 9600 9680 9640 9720
rect 9680 9680 9720 9720
rect 9760 9680 9800 9720
rect 9840 9680 9890 9720
rect 9930 9680 9970 9720
rect 10010 9680 10050 9720
rect 10090 9680 10130 9720
rect 10170 9680 10210 9720
rect 10250 9680 10290 9720
rect 10330 9680 10370 9720
rect 10410 9680 10450 9720
rect 10490 9680 10530 9720
rect 10570 9680 10610 9720
rect 10650 9680 10690 9720
rect 10730 9680 10770 9720
rect 10810 9680 10850 9720
rect 10890 9680 10930 9720
rect 10970 9680 11010 9720
rect 11050 9680 11090 9720
rect 11130 9680 11170 9720
rect 11210 9680 11250 9720
rect 11290 9680 11330 9720
rect 11370 9680 11410 9720
rect 11450 9680 11490 9720
rect 11530 9680 11570 9720
rect 11610 9680 11650 9720
rect 11690 9680 11730 9720
rect 11770 9680 11810 9720
rect 11850 9680 11890 9720
rect 11930 9680 11970 9720
rect 12010 9680 12050 9720
rect 12090 9680 12130 9720
rect 12170 9680 12210 9720
rect 12250 9680 12290 9720
rect 12330 9680 12370 9720
rect 12410 9680 12450 9720
rect 12490 9680 12530 9720
rect 12570 9680 12610 9720
rect 12650 9680 12690 9720
rect 12730 9680 12770 9720
rect 12810 9680 12850 9720
rect 12890 9680 12930 9720
rect 12970 9680 13010 9720
rect 13050 9680 13090 9720
rect 13130 9680 13170 9720
rect 13210 9680 13250 9720
rect 13290 9680 13330 9720
rect 13370 9680 13410 9720
rect 13450 9680 13490 9720
rect 13530 9680 13570 9720
rect 13610 9680 13650 9720
rect 13690 9680 13730 9720
rect 13770 9680 13810 9720
rect 13850 9680 13890 9720
rect 13930 9680 13970 9720
rect 14010 9680 14050 9720
rect 14090 9680 14130 9720
rect 14170 9680 14210 9720
rect 14250 9680 14290 9720
rect 14330 9680 14370 9720
rect 14410 9680 14450 9720
rect 14490 9680 14530 9720
rect 14570 9680 14610 9720
rect 14650 9680 14690 9720
rect 14730 9680 14770 9720
rect 14810 9680 14850 9720
rect 14890 9680 14930 9720
rect 14970 9680 15010 9720
rect 15050 9680 15090 9720
rect 15130 9680 15170 9720
rect 15210 9680 15250 9720
rect 15290 9680 15330 9720
rect 15370 9680 15410 9720
rect 15450 9680 15490 9720
rect 15530 9680 15570 9720
rect 15610 9680 15650 9720
rect 15690 9680 15730 9720
rect 15770 9680 15810 9720
rect 15850 9680 15890 9720
rect 15930 9680 15970 9720
rect 16010 9680 16050 9720
rect 16090 9680 16130 9720
rect 16170 9680 16210 9720
rect 16250 9680 16290 9720
rect 16330 9680 16370 9720
rect 16410 9680 16450 9720
rect 16490 9680 16530 9720
rect 16570 9680 16610 9720
rect 16650 9680 16690 9720
rect 16730 9680 16770 9720
rect 16810 9680 16850 9720
rect 16890 9680 16930 9720
rect 16970 9680 17010 9720
rect 17050 9680 17090 9720
rect 17130 9680 17170 9720
rect 17210 9680 17250 9720
rect 17290 9680 17330 9720
rect 17370 9680 17410 9720
rect 17450 9680 17490 9720
rect 17530 9680 17570 9720
rect 17610 9680 17650 9720
rect 17690 9680 17730 9720
rect 17770 9680 17810 9720
rect 17850 9680 17890 9720
rect 17930 9680 17970 9720
rect 18010 9680 18050 9720
rect 18090 9680 18130 9720
rect 18170 9680 18210 9720
rect 18250 9680 18290 9720
rect 18330 9680 18370 9720
rect 18410 9680 18450 9720
rect 18490 9680 18530 9720
rect 18570 9680 18610 9720
rect 18650 9680 18690 9720
rect 18730 9680 18770 9720
rect 18810 9680 18850 9720
rect 18890 9680 18930 9720
rect 18970 9680 19010 9720
rect 19050 9680 19090 9720
rect 19130 9680 19170 9720
rect 19210 9680 19250 9720
rect 19290 9680 19330 9720
rect 19370 9680 19410 9720
rect 19450 9680 19490 9720
rect 19530 9680 19570 9720
rect 19610 9680 19650 9720
rect 19690 9680 19730 9720
rect 19770 9680 19810 9720
rect 19850 9680 19890 9720
rect 19930 9680 19970 9720
rect 20010 9680 20050 9720
rect 20090 9680 20130 9720
rect 20170 9680 20210 9720
rect 20250 9680 20290 9720
rect 20330 9680 20370 9720
rect 20410 9680 20450 9720
rect 20490 9680 20530 9720
rect 20570 9680 20610 9720
rect 20650 9680 20690 9720
rect 20730 9680 20770 9720
rect 20810 9680 20850 9720
rect 20890 9680 20930 9720
rect 20970 9680 21010 9720
rect 21050 9680 21160 9720
rect 8470 9650 21160 9680
rect 7280 9630 21160 9650
rect 7280 9590 7740 9630
rect 7780 9590 7820 9630
rect 7860 9590 7900 9630
rect 7940 9590 7980 9630
rect 8020 9590 8060 9630
rect 8100 9590 8140 9630
rect 8180 9590 8220 9630
rect 8260 9590 8300 9630
rect 8340 9590 8380 9630
rect 8420 9590 8460 9630
rect 8500 9610 21160 9630
rect 8500 9590 8880 9610
rect 7280 8800 8880 9590
rect 9690 8800 9910 9610
rect 10720 8800 10940 9610
rect 11750 8800 11970 9610
rect 12780 8800 12980 9610
rect 13790 8800 14010 9610
rect 14820 8800 15040 9610
rect 15850 8800 16070 9610
rect 16880 8800 17080 9610
rect 17890 8800 18110 9610
rect 18920 8800 19120 9610
rect 19930 8800 20150 9610
rect 21110 8800 21160 9610
rect 21570 8940 21640 10340
rect 21970 8940 22040 12640
rect 22400 8940 22470 14960
rect 21550 8920 21660 8940
rect 21550 8850 21570 8920
rect 21640 8850 21660 8920
rect 21550 8830 21660 8850
rect 21950 8920 22060 8940
rect 21950 8850 21970 8920
rect 22040 8850 22060 8920
rect 21950 8830 22060 8850
rect 22380 8920 22490 8940
rect 22380 8850 22400 8920
rect 22470 8850 22490 8920
rect 22380 8830 22490 8850
rect 7280 8750 21160 8800
rect 22550 8640 22660 8660
rect 13190 8630 22570 8640
rect 13190 8580 13220 8630
rect 13270 8580 22570 8630
rect 13190 8570 22570 8580
rect 22640 8570 22660 8640
rect 22550 8550 22660 8570
rect 13390 8490 13600 8510
rect 13390 8420 13430 8490
rect 13560 8420 13600 8490
rect 13190 8230 13300 8420
rect 13390 8400 13600 8420
rect 22760 8370 22860 18290
rect 17020 8360 22860 8370
rect 17020 8310 17050 8360
rect 17100 8310 22860 8360
rect 17020 8300 22860 8310
rect 12100 6990 12160 7000
rect 9870 6980 17060 6990
rect 9870 6930 9900 6980
rect 9960 6930 10120 6980
rect 10180 6930 10340 6980
rect 10400 6930 10560 6980
rect 10620 6930 10780 6980
rect 10840 6930 11000 6980
rect 11060 6930 11220 6980
rect 11280 6930 11440 6980
rect 11500 6930 11660 6980
rect 11720 6930 11880 6980
rect 11940 6930 12100 6980
rect 12160 6930 12320 6980
rect 12380 6930 12540 6980
rect 12600 6930 12760 6980
rect 12820 6930 12980 6980
rect 13040 6930 13200 6980
rect 13260 6930 13670 6980
rect 13730 6930 13890 6980
rect 13950 6930 14110 6980
rect 14170 6930 14330 6980
rect 14390 6930 14550 6980
rect 14610 6930 14770 6980
rect 14830 6930 14990 6980
rect 15050 6930 15210 6980
rect 15270 6930 15430 6980
rect 15490 6930 15650 6980
rect 15710 6930 15870 6980
rect 15930 6930 16090 6980
rect 16150 6930 16310 6980
rect 16370 6930 16530 6980
rect 16590 6930 16750 6980
rect 16810 6930 16970 6980
rect 17030 6930 17060 6980
rect 9870 6870 17060 6930
rect 9870 6060 9930 6870
rect 11200 6060 11430 6870
rect 12240 6060 12460 6870
rect 13270 6060 13660 6870
rect 14930 6060 15160 6870
rect 15970 6060 16190 6870
rect 17000 6060 17060 6870
rect 9870 5990 17060 6060
rect 9870 5960 13630 5990
rect 13600 5940 13630 5960
rect 13690 5940 13850 5990
rect 13910 5940 14070 5990
rect 14130 5940 14290 5990
rect 14350 5940 14510 5990
rect 14570 5940 14730 5990
rect 14790 5940 14950 5990
rect 15010 5940 15170 5990
rect 15230 5940 15390 5990
rect 15450 5940 15610 5990
rect 15670 5940 15830 5990
rect 15890 5940 16050 5990
rect 16110 5940 16270 5990
rect 16330 5940 16490 5990
rect 16550 5940 16710 5990
rect 16770 5940 16930 5990
rect 16990 5940 17060 5990
rect 13600 5930 17060 5940
rect 15830 5920 15890 5930
rect 13340 5880 13550 5900
rect 9870 5870 13170 5880
rect 9870 5830 9930 5870
rect 9970 5830 10010 5870
rect 10050 5830 10090 5870
rect 10130 5830 10170 5870
rect 10210 5830 10250 5870
rect 10290 5830 10330 5870
rect 10370 5830 10410 5870
rect 10450 5830 10490 5870
rect 10530 5830 10610 5870
rect 10650 5830 10690 5870
rect 10730 5830 10770 5870
rect 10810 5830 10850 5870
rect 10890 5830 10930 5870
rect 10970 5830 11010 5870
rect 11050 5830 11090 5870
rect 11130 5830 11170 5870
rect 11210 5830 11250 5870
rect 11290 5830 11370 5870
rect 11410 5830 11450 5870
rect 11490 5830 11530 5870
rect 11570 5830 11610 5870
rect 11650 5830 11690 5870
rect 11730 5830 11770 5870
rect 11810 5830 11850 5870
rect 11890 5830 11930 5870
rect 11970 5830 12010 5870
rect 12050 5830 12130 5870
rect 12170 5830 12210 5870
rect 12250 5830 12290 5870
rect 12330 5830 12370 5870
rect 12410 5830 12450 5870
rect 12490 5830 12530 5870
rect 12570 5830 12610 5870
rect 12650 5830 12690 5870
rect 12730 5830 12770 5870
rect 12810 5830 12850 5870
rect 12890 5830 12930 5870
rect 12970 5830 13010 5870
rect 13050 5830 13090 5870
rect 13130 5830 13170 5870
rect 9870 5820 13170 5830
rect 13340 5820 13380 5880
rect 13510 5820 13550 5880
rect 13340 5800 13550 5820
rect 13400 4520 13490 5800
rect 13340 4500 13550 4520
rect 13340 4440 13380 4500
rect 13510 4440 13550 4500
rect 23070 4480 23140 22620
rect 23250 8640 23360 8660
rect 23430 8640 23510 24880
rect 23250 8570 23270 8640
rect 23340 8570 23510 8640
rect 23250 8550 23360 8570
rect 13340 4420 13550 4440
rect 16920 4470 23140 4480
rect 16920 4420 16950 4470
rect 17000 4420 23140 4470
rect 16920 4410 23140 4420
rect 13340 4340 13550 4360
rect 13340 4280 13380 4340
rect 13510 4280 13550 4340
rect 13340 4260 13550 4280
rect 21950 4310 22060 4330
rect 21950 4240 21970 4310
rect 22040 4240 22060 4310
rect 21950 4220 22060 4240
rect 22380 4310 22490 4330
rect 22380 4240 22400 4310
rect 22470 4240 22490 4310
rect 22380 4220 22490 4240
rect 19180 4170 19330 4200
rect 9840 4140 9940 4160
rect 9840 4070 9850 4140
rect 9930 4070 9940 4140
rect 13160 4150 19200 4170
rect 13160 4090 13180 4150
rect 13250 4090 19200 4150
rect 13160 4070 19200 4090
rect 19310 4070 19330 4170
rect 9840 4050 9940 4070
rect 19180 4040 19330 4070
rect 200 3990 600 4010
rect 200 3880 230 3990
rect 570 3980 600 3990
rect 570 3960 13270 3980
rect 570 3900 13180 3960
rect 13250 3900 13270 3960
rect 570 3880 13270 3900
rect 200 3860 600 3880
rect 21970 3250 22040 4220
rect 16920 3240 22040 3250
rect 16920 3190 16950 3240
rect 17000 3190 22040 3240
rect 16920 3180 22040 3190
rect 13280 3080 13490 3100
rect 13280 3020 13320 3080
rect 13450 3020 13490 3080
rect 13280 3000 13490 3020
rect 13600 3000 17060 3010
rect 13600 2950 13630 3000
rect 13690 2950 13850 3000
rect 13910 2950 14070 3000
rect 14130 2950 14290 3000
rect 14350 2950 14510 3000
rect 14570 2950 14730 3000
rect 14790 2950 14950 3000
rect 15010 2950 15170 3000
rect 15230 2950 15390 3000
rect 15450 2950 15610 3000
rect 15670 2950 15830 3000
rect 15890 2950 16050 3000
rect 16110 2950 16270 3000
rect 16330 2950 16490 3000
rect 16550 2950 16710 3000
rect 16770 2950 17060 3000
rect 13600 2940 17060 2950
rect 9850 2840 17060 2940
rect 9850 2030 9910 2840
rect 11130 2030 11350 2840
rect 12160 2030 12370 2840
rect 13180 2030 13570 2840
rect 14950 2030 15170 2840
rect 15980 2030 16190 2840
rect 17000 2030 17060 2840
rect 9850 1920 17060 2030
rect 9850 1870 9890 1920
rect 9950 1870 10110 1920
rect 10170 1870 10330 1920
rect 10390 1870 10550 1920
rect 10610 1870 10770 1920
rect 10830 1870 10990 1920
rect 11050 1870 11210 1920
rect 11270 1870 11430 1920
rect 11490 1870 11650 1920
rect 11710 1870 11870 1920
rect 11930 1870 12090 1920
rect 12150 1870 12310 1920
rect 12370 1870 12530 1920
rect 12590 1870 12750 1920
rect 12810 1870 12970 1920
rect 13030 1870 13630 1920
rect 13690 1870 13850 1920
rect 13910 1870 14070 1920
rect 14130 1870 14290 1920
rect 14350 1870 14510 1920
rect 14570 1870 14730 1920
rect 14790 1870 14950 1920
rect 15010 1870 15170 1920
rect 15230 1870 15390 1920
rect 15450 1870 15610 1920
rect 15670 1870 15830 1920
rect 15890 1870 16050 1920
rect 16110 1870 16270 1920
rect 16330 1870 16490 1920
rect 16550 1870 16710 1920
rect 16770 1870 17060 1920
rect 9850 1860 17060 1870
rect 13180 1680 13610 1690
rect 13180 1630 13210 1680
rect 13260 1630 13610 1680
rect 13180 1620 13610 1630
rect 13320 600 13530 620
rect 13320 530 13360 600
rect 13490 530 13530 600
rect 13320 510 13530 530
rect 13560 420 13610 1620
rect 22400 1430 22470 4220
rect 25790 2780 27600 2810
rect 23110 2720 24290 2770
rect 23110 2710 24220 2720
rect 23110 2080 23170 2710
rect 23980 2660 24220 2710
rect 24280 2660 24290 2720
rect 23980 2620 24290 2660
rect 23980 2560 24220 2620
rect 24280 2560 24290 2620
rect 23980 2520 24290 2560
rect 23980 2460 24220 2520
rect 24280 2460 24290 2520
rect 23980 2420 24290 2460
rect 23980 2360 24220 2420
rect 24280 2360 24290 2420
rect 23980 2320 24290 2360
rect 23980 2260 24220 2320
rect 24280 2260 24290 2320
rect 23980 2220 24290 2260
rect 23980 2160 24220 2220
rect 24280 2160 24290 2220
rect 23980 2120 24290 2160
rect 23980 2080 24220 2120
rect 23110 2060 24220 2080
rect 24280 2060 24290 2120
rect 25710 2760 27230 2780
rect 25710 2720 25720 2760
rect 25770 2720 27230 2760
rect 25710 2640 27230 2720
rect 25710 2600 25720 2640
rect 25770 2600 27230 2640
rect 25710 2520 27230 2600
rect 25710 2480 25720 2520
rect 25770 2480 27230 2520
rect 25710 2400 27230 2480
rect 25710 2360 25720 2400
rect 25770 2360 27230 2400
rect 25710 2280 27230 2360
rect 25710 2240 25720 2280
rect 25770 2240 27230 2280
rect 25710 2160 27230 2240
rect 25710 2120 25720 2160
rect 25770 2130 27230 2160
rect 27570 2130 27600 2780
rect 25770 2120 27600 2130
rect 25710 2100 27600 2120
rect 23110 2030 24290 2060
rect 25810 2030 26090 2100
rect 25470 1970 26090 2030
rect 25470 1910 25480 1970
rect 25540 1910 26090 1970
rect 25470 1860 26090 1910
rect 17030 1420 22470 1430
rect 17030 1370 17060 1420
rect 17110 1370 22470 1420
rect 17030 1360 22470 1370
rect 21550 420 21660 440
rect 13560 350 21570 420
rect 21640 350 21660 420
rect 21550 330 21660 350
<< via1 >>
rect 2120 43410 2950 44100
rect 21730 43410 22580 44100
rect 22980 43410 23830 44100
rect 21830 43280 21890 43350
rect 21930 43280 21990 43350
rect 22030 43280 22090 43350
rect 22130 43280 22190 43350
rect 22230 43280 22290 43350
rect 22330 43280 22390 43350
rect 22430 43280 22490 43350
rect 22530 43280 22590 43350
rect 22630 43280 22690 43350
rect 22730 43280 22790 43350
rect 22830 43280 22890 43350
rect 22930 43280 22990 43350
rect 23030 43280 23090 43350
rect 23130 43280 23190 43350
rect 23230 43280 23290 43350
rect 23330 43280 23390 43350
rect 23430 43280 23490 43350
rect 23530 43280 23590 43350
rect 15690 43050 15770 43180
rect 22340 43090 22400 43150
rect 3430 42310 4280 43000
rect 3079 41680 3179 41690
rect 3079 41640 3089 41680
rect 3089 41640 3169 41680
rect 3169 41640 3179 41680
rect 3079 41630 3179 41640
rect 3179 41460 3239 41520
rect 5509 40860 5569 40920
rect 6009 41910 6069 41970
rect 6119 41910 6179 41970
rect 6229 41910 6289 41970
rect 6339 41910 6399 41970
rect 6449 41910 6509 41970
rect 6559 41910 6619 41970
rect 6669 41910 6729 41970
rect 6779 41910 6839 41970
rect 6889 41910 6949 41970
rect 6999 41910 7059 41970
rect 7109 41910 7169 41970
rect 7219 41910 7279 41970
rect 7329 41910 7389 41970
rect 7439 41910 7499 41970
rect 7549 41910 7609 41970
rect 7659 41910 7719 41970
rect 7769 41910 7829 41970
rect 7879 41910 7939 41970
rect 7989 41910 8049 41970
rect 8099 41910 8159 41970
rect 8209 41910 8269 41970
rect 8319 41910 8379 41970
rect 8429 41910 8489 41970
rect 8539 41910 8599 41970
rect 8649 41910 8709 41970
rect 8759 41910 8819 41970
rect 8869 41910 8929 41970
rect 8979 41910 9039 41970
rect 9089 41910 9149 41970
rect 9199 41910 9259 41970
rect 9309 41910 9369 41970
rect 9419 41910 9479 41970
rect 9529 41910 9589 41970
rect 9639 41910 9699 41970
rect 9749 41910 9809 41970
rect 9859 41910 9919 41970
rect 22070 42070 22130 42130
rect 23640 41810 23720 41870
rect 22450 41270 22510 41330
rect 21620 41090 21680 41160
rect 21720 41090 21780 41160
rect 21830 41090 21890 41160
rect 21930 41090 21990 41160
rect 22030 41090 22090 41160
rect 22130 41090 22190 41160
rect 22230 41090 22290 41160
rect 22330 41090 22390 41160
rect 22430 41090 22490 41160
rect 22530 41090 22590 41160
rect 22630 41090 22690 41160
rect 22730 41090 22790 41160
rect 22830 41090 22890 41160
rect 22930 41090 22990 41160
rect 23030 41090 23090 41160
rect 23130 41090 23190 41160
rect 23230 41090 23290 41160
rect 23330 41090 23390 41160
rect 23430 41090 23490 41160
rect 23530 41090 23590 41160
rect 6409 40590 6469 40650
rect 6519 40590 6579 40650
rect 6629 40590 6689 40650
rect 6739 40590 6799 40650
rect 6849 40590 6909 40650
rect 6959 40590 7019 40650
rect 7069 40590 7129 40650
rect 7179 40590 7239 40650
rect 7289 40590 7349 40650
rect 7399 40590 7459 40650
rect 7509 40590 7569 40650
rect 7619 40590 7679 40650
rect 7729 40590 7789 40650
rect 7839 40590 7899 40650
rect 7949 40590 8009 40650
rect 8059 40590 8119 40650
rect 8169 40590 8229 40650
rect 8279 40590 8339 40650
rect 8389 40590 8449 40650
rect 8499 40590 8559 40650
rect 8609 40590 8669 40650
rect 8719 40590 8779 40650
rect 8829 40590 8889 40650
rect 8939 40590 8999 40650
rect 9049 40590 9109 40650
rect 9159 40590 9219 40650
rect 9269 40590 9329 40650
rect 9379 40590 9439 40650
rect 9489 40590 9549 40650
rect 9599 40590 9659 40650
rect 9709 40590 9769 40650
rect 9819 40590 9879 40650
rect 21610 40340 22250 41020
rect 22440 40340 23080 41020
rect 23260 40340 23900 41020
rect 10060 39880 10900 40000
rect 3149 39500 3209 39560
rect 2130 38620 3170 39430
rect 3380 38620 4420 39430
rect 4630 38620 5670 39430
rect 5880 38620 6920 39430
rect 7130 38620 8170 39430
rect 8380 38620 9850 39430
rect 25330 38430 25400 38500
rect 25840 38430 25910 38500
rect 2120 37240 3860 38050
rect 4070 37240 5110 38050
rect 5320 37240 6360 38050
rect 6570 37240 7610 38050
rect 7820 37240 8860 38050
rect 9070 37240 9820 38050
rect 10080 37240 10880 38050
rect 12970 36400 13760 37200
rect 13970 36400 14760 37200
rect 4560 34930 4620 35000
rect 2120 32670 2950 33360
rect 3150 32670 3980 33360
rect 4180 32670 5010 33360
rect 5210 32670 6040 33360
rect 6240 32670 7070 33360
rect 7270 32670 8100 33360
rect 8300 32670 9130 33360
rect 9330 32670 10870 33360
rect 2120 31790 2950 32480
rect 3150 31790 3980 32480
rect 4180 31790 5010 32480
rect 5210 31790 6040 32480
rect 6240 31790 7070 32480
rect 7270 31790 8100 32480
rect 8300 31790 9130 32480
rect 9330 31790 10160 32480
rect 10360 31790 11190 32480
rect 2960 30680 3020 30740
rect 2120 28310 2950 29000
rect 3150 28310 3980 29000
rect 4180 28310 5010 29000
rect 5210 28310 6040 29000
rect 6240 28310 7070 29000
rect 7270 28310 8100 29000
rect 8300 28310 9130 29000
rect 9330 28310 10160 29000
rect 10360 28310 11190 29000
rect 5380 27990 5480 28100
rect 5610 27710 5710 27820
rect 6300 25500 6360 25560
rect 15570 35570 15640 35630
rect 15790 35570 15900 35630
rect 16450 35430 16510 35490
rect 17240 35240 17310 35310
rect 20730 36090 20790 36170
rect 20730 35830 20790 35910
rect 18270 35230 18340 35300
rect 18310 34540 18370 34620
rect 19750 34750 19810 34810
rect 20920 34900 20980 34960
rect 22200 35240 22270 35310
rect 23520 35170 23590 35240
rect 20760 34450 20820 34530
rect 19580 34350 19640 34430
rect 23240 34470 23300 34550
rect 24710 34750 24770 34810
rect 24950 34300 25010 34380
rect 22440 33250 23080 34060
rect 15650 32250 15710 32310
rect 14400 31950 14510 32010
rect 15590 31940 15650 32020
rect 15400 30210 15470 30280
rect 16450 31390 16510 31450
rect 17240 31230 17310 31300
rect 18540 31080 18610 31150
rect 18240 30400 18310 30480
rect 20010 30690 20070 30750
rect 20740 30760 20800 30840
rect 20980 30840 21040 30900
rect 22260 31230 22330 31300
rect 23570 31080 23640 31150
rect 20560 30380 20620 30460
rect 20740 30380 20800 30460
rect 23260 30400 23320 30480
rect 24970 30680 25030 30740
rect 22440 29170 23080 29980
rect 12720 28510 12820 28620
rect 12710 28160 12810 28270
rect 7370 26670 8200 27360
rect 8400 26670 9230 27360
rect 9430 26670 10260 27360
rect 10460 26670 11290 27360
rect 11490 26670 12320 27360
rect 12520 26670 13350 27360
rect 13550 26670 14380 27360
rect 14580 26670 15410 27360
rect 15610 26670 16440 27360
rect 16640 26670 17470 27360
rect 17670 26670 18500 27360
rect 18700 26670 19530 27360
rect 19760 26670 20590 27360
rect 8080 24800 8140 24870
rect 7570 24710 7630 24770
rect 10410 24790 10480 24850
rect 11410 24790 11480 24850
rect 8200 24670 8260 24730
rect 9090 24380 9160 24440
rect 19560 23380 20370 24190
rect 9090 23080 9160 23140
rect 10410 22720 10480 22780
rect 11410 22720 11480 22780
rect 9220 22640 9280 22700
rect 12730 20350 12800 20410
rect 17670 20090 18500 20890
rect 7110 19410 7170 19470
rect 6960 18620 7020 18680
rect 7230 18360 7290 18420
rect 9220 18270 9280 18330
rect 10410 18200 10480 18260
rect 9470 18040 9540 18100
rect 9090 17900 9160 17960
rect 19560 16790 20370 17600
rect 10920 15720 11750 16410
rect 11950 15720 12780 16410
rect 12980 15720 13810 16410
rect 14040 15720 14870 16410
rect 15070 15720 15900 16410
rect 16100 15720 16930 16410
rect 17160 15720 17990 16410
rect 18190 15720 19020 16410
rect 19220 15720 20050 16410
rect 20280 15720 21110 16410
rect 7430 15230 7500 15290
rect 9750 15050 9810 15110
rect 10280 14960 10350 15020
rect 8430 14200 8500 14260
rect 9910 13430 10720 14240
rect 10940 13430 11750 14240
rect 11970 13430 12780 14240
rect 12980 13430 13790 14240
rect 7700 12650 7760 12710
rect 7590 12540 7650 12600
rect 9670 13090 9740 13150
rect 11280 12550 11350 12610
rect 9750 12470 9820 12530
rect 14040 11170 14870 11860
rect 15070 11170 15900 11860
rect 16100 11170 16930 11860
rect 17160 11170 17990 11860
rect 18190 11170 19020 11860
rect 19220 11170 20050 11860
rect 20280 11170 21110 11860
rect 7610 10890 7670 10950
rect 7850 10790 7910 10850
rect 9650 10780 9720 10840
rect 11290 10470 11360 10530
rect 9790 10350 9860 10410
rect 12290 10440 12360 10500
rect 8880 8800 9690 9610
rect 9910 8800 10720 9610
rect 10940 8800 11750 9610
rect 11970 8800 12780 9610
rect 12980 8800 13790 9610
rect 14010 8800 14820 9610
rect 15040 8800 15850 9610
rect 16070 8800 16880 9610
rect 17080 8800 17890 9610
rect 18110 8800 18920 9610
rect 19120 8800 19930 9610
rect 20150 8800 21110 9610
rect 21570 8850 21640 8920
rect 21970 8850 22040 8920
rect 22400 8850 22470 8920
rect 22570 8570 22640 8640
rect 13430 8420 13560 8490
rect 9930 6060 11200 6870
rect 11430 6060 12240 6870
rect 12460 6060 13270 6870
rect 13660 6060 14930 6870
rect 15160 6060 15970 6870
rect 16190 6060 17000 6870
rect 13380 5820 13510 5880
rect 13380 4440 13510 4500
rect 23270 8570 23340 8640
rect 13380 4280 13510 4340
rect 21970 4240 22040 4310
rect 22400 4240 22470 4310
rect 9850 4070 9930 4140
rect 19200 4070 19310 4170
rect 230 3880 570 3990
rect 13320 3020 13450 3080
rect 9910 2030 11130 2840
rect 11350 2030 12160 2840
rect 12370 2030 13180 2840
rect 13570 2030 14950 2840
rect 15170 2030 15980 2840
rect 16190 2030 17000 2840
rect 13360 530 13490 600
rect 23170 2080 23980 2710
rect 27230 2130 27570 2780
rect 21570 350 21640 420
<< metal2 >>
rect 24500 44560 24620 44580
rect 11570 44430 24520 44560
rect 24600 44430 24620 44560
rect 2070 44100 3000 44160
rect 2070 43410 2120 44100
rect 2950 43410 3000 44100
rect 2070 43360 3000 43410
rect 3380 43000 4330 43060
rect 3380 42310 3430 43000
rect 4280 42310 4330 43000
rect 3380 42260 4330 42310
rect 5949 41970 9979 41980
rect 5949 41910 6009 41970
rect 6069 41910 6119 41970
rect 6179 41910 6229 41970
rect 6289 41910 6339 41970
rect 6399 41910 6449 41970
rect 6509 41910 6559 41970
rect 6619 41910 6669 41970
rect 6729 41910 6779 41970
rect 6839 41910 6889 41970
rect 6949 41910 6999 41970
rect 7059 41910 7109 41970
rect 7169 41910 7219 41970
rect 7279 41910 7329 41970
rect 7389 41910 7439 41970
rect 7499 41910 7549 41970
rect 7609 41910 7659 41970
rect 7719 41910 7769 41970
rect 7829 41910 7879 41970
rect 7939 41910 7989 41970
rect 8049 41910 8099 41970
rect 8159 41910 8209 41970
rect 8269 41910 8319 41970
rect 8379 41910 8429 41970
rect 8489 41910 8539 41970
rect 8599 41910 8649 41970
rect 8709 41910 8759 41970
rect 8819 41910 8869 41970
rect 8929 41910 8979 41970
rect 9039 41910 9089 41970
rect 9149 41910 9199 41970
rect 9259 41910 9309 41970
rect 9369 41910 9419 41970
rect 9479 41910 9529 41970
rect 9589 41910 9639 41970
rect 9699 41910 9749 41970
rect 9809 41910 9859 41970
rect 9919 41910 9979 41970
rect 5949 41900 9979 41910
rect 3049 41690 3209 41700
rect 3049 41630 3079 41690
rect 3179 41630 3209 41690
rect 3049 41620 3209 41630
rect 3089 40840 3129 41620
rect 3159 41520 3259 41530
rect 3159 41460 3179 41520
rect 3239 41460 3259 41520
rect 3159 41450 3259 41460
rect 3179 40910 3219 41450
rect 5489 40920 5589 40930
rect 5489 40910 5509 40920
rect 3179 40870 5509 40910
rect 5489 40860 5509 40870
rect 5569 40860 5589 40920
rect 5489 40850 5589 40860
rect 3089 40800 3199 40840
rect 3159 39570 3199 40800
rect 6129 40790 6169 41900
rect 6129 40770 9879 40790
rect 6129 40740 9880 40770
rect 6350 40660 9880 40740
rect 6349 40650 9969 40660
rect 6349 40590 6409 40650
rect 6469 40590 6519 40650
rect 6579 40590 6629 40650
rect 6689 40590 6739 40650
rect 6799 40590 6849 40650
rect 6909 40590 6959 40650
rect 7019 40590 7069 40650
rect 7129 40590 7179 40650
rect 7239 40590 7289 40650
rect 7349 40590 7399 40650
rect 7459 40590 7509 40650
rect 7569 40590 7619 40650
rect 7679 40590 7729 40650
rect 7789 40590 7839 40650
rect 7899 40590 7949 40650
rect 8009 40590 8059 40650
rect 8119 40590 8169 40650
rect 8229 40590 8279 40650
rect 8339 40590 8389 40650
rect 8449 40590 8499 40650
rect 8559 40590 8609 40650
rect 8669 40590 8719 40650
rect 8779 40590 8829 40650
rect 8889 40590 8939 40650
rect 8999 40590 9049 40650
rect 9109 40590 9159 40650
rect 9219 40590 9269 40650
rect 9329 40590 9379 40650
rect 9439 40590 9489 40650
rect 9549 40590 9599 40650
rect 9659 40590 9709 40650
rect 9769 40590 9819 40650
rect 9879 40590 9969 40650
rect 6349 40580 9969 40590
rect 10030 40000 10930 40020
rect 10030 39880 10060 40000
rect 10900 39880 10930 40000
rect 10030 39860 10930 39880
rect 3139 39560 3219 39570
rect 3139 39500 3149 39560
rect 3209 39500 3219 39560
rect 3139 39490 3219 39500
rect 2070 39430 3220 39490
rect 2070 38620 2130 39430
rect 3170 38620 3220 39430
rect 2070 38560 3220 38620
rect 3320 39430 4470 39490
rect 3320 38620 3380 39430
rect 4420 38620 4470 39430
rect 3320 38560 4470 38620
rect 4570 39430 5720 39490
rect 4570 38620 4630 39430
rect 5670 38620 5720 39430
rect 4570 38560 5720 38620
rect 5820 39430 6970 39490
rect 5820 38620 5880 39430
rect 6920 38620 6970 39430
rect 5820 38560 6970 38620
rect 7070 39430 8220 39490
rect 7070 38620 7130 39430
rect 8170 38620 8220 39430
rect 7070 38560 8220 38620
rect 8320 39430 9900 39490
rect 8320 38620 8380 39430
rect 9850 38620 9900 39430
rect 8320 38560 9900 38620
rect 2070 38050 3910 38110
rect 2070 37240 2120 38050
rect 3860 37240 3910 38050
rect 2070 37180 3910 37240
rect 4010 38050 5160 38110
rect 4010 37240 4070 38050
rect 5110 37240 5160 38050
rect 4010 37180 5160 37240
rect 5260 38050 6410 38110
rect 5260 37240 5320 38050
rect 6360 37240 6410 38050
rect 5260 37180 6410 37240
rect 6510 38050 7660 38110
rect 6510 37240 6570 38050
rect 7610 37240 7660 38050
rect 6510 37180 7660 37240
rect 7760 38050 8910 38110
rect 7760 37240 7820 38050
rect 8860 37240 8910 38050
rect 7760 37180 8910 37240
rect 9010 38050 9870 38110
rect 9010 37240 9070 38050
rect 9820 37240 9870 38050
rect 9010 37180 9870 37240
rect 10030 38050 10930 38110
rect 10030 37240 10080 38050
rect 10880 37240 10930 38050
rect 10030 37180 10930 37240
rect 11570 35720 11700 44430
rect 24500 44410 24620 44430
rect 25600 44560 25720 44580
rect 25600 44430 25620 44560
rect 25700 44430 25720 44560
rect 25600 44410 25720 44430
rect 26150 44560 26270 44580
rect 26150 44430 26170 44560
rect 26250 44430 26270 44560
rect 26150 44410 26270 44430
rect 21680 44100 22630 44160
rect 21680 43410 21730 44100
rect 22580 43410 22630 44100
rect 21680 43360 22630 43410
rect 22930 44100 23880 44160
rect 22930 43410 22980 44100
rect 23830 43410 23880 44100
rect 22930 43360 23880 43410
rect 21790 43350 23630 43360
rect 21790 43280 21830 43350
rect 21890 43280 21930 43350
rect 21990 43280 22030 43350
rect 22090 43280 22130 43350
rect 22190 43280 22230 43350
rect 22290 43280 22330 43350
rect 22390 43280 22430 43350
rect 22490 43280 22530 43350
rect 22590 43280 22630 43350
rect 22690 43280 22730 43350
rect 22790 43280 22830 43350
rect 22890 43280 22930 43350
rect 22990 43280 23030 43350
rect 23090 43280 23130 43350
rect 23190 43280 23230 43350
rect 23290 43280 23330 43350
rect 23390 43280 23430 43350
rect 23490 43280 23530 43350
rect 23590 43280 23630 43350
rect 21790 43270 23630 43280
rect 15670 43180 15790 43200
rect 15670 43050 15690 43180
rect 15770 43050 15790 43180
rect 22320 43150 22420 43170
rect 22320 43090 22340 43150
rect 22400 43090 22420 43150
rect 22320 43070 22420 43090
rect 15670 43030 15790 43050
rect 22050 42130 22150 42140
rect 22050 42070 22070 42130
rect 22130 42070 22150 42130
rect 22050 41590 22150 42070
rect 21290 41500 22150 41590
rect 21290 38510 21390 41500
rect 22350 41180 22390 43070
rect 22460 41350 22500 43270
rect 23620 41870 23740 41890
rect 23620 41810 23640 41870
rect 23720 41810 23740 41870
rect 23620 41790 23740 41810
rect 22430 41330 22530 41350
rect 22430 41270 22450 41330
rect 22510 41270 22530 41330
rect 22430 41250 22530 41270
rect 21590 41160 23630 41180
rect 21590 41090 21620 41160
rect 21680 41090 21720 41160
rect 21780 41090 21830 41160
rect 21890 41090 21930 41160
rect 21990 41090 22030 41160
rect 22090 41090 22130 41160
rect 22190 41090 22230 41160
rect 22290 41090 22330 41160
rect 22390 41090 22430 41160
rect 22490 41090 22530 41160
rect 22590 41090 22630 41160
rect 22690 41090 22730 41160
rect 22790 41090 22830 41160
rect 22890 41090 22930 41160
rect 22990 41090 23030 41160
rect 23090 41090 23130 41160
rect 23190 41090 23230 41160
rect 23290 41090 23330 41160
rect 23390 41090 23430 41160
rect 23490 41090 23530 41160
rect 23590 41090 23630 41160
rect 21590 41080 23630 41090
rect 21560 41020 22300 41080
rect 21560 40340 21610 41020
rect 22250 40340 22300 41020
rect 21560 40290 22300 40340
rect 22390 41020 23130 41080
rect 22390 40340 22440 41020
rect 23080 40340 23130 41020
rect 22390 40290 23130 40340
rect 23210 41020 23950 41080
rect 23210 40340 23260 41020
rect 23900 40340 23950 41020
rect 23210 40290 23950 40340
rect 25320 38510 25410 38520
rect 1890 35610 11700 35720
rect 11930 38500 25410 38510
rect 11930 38430 25330 38500
rect 25400 38430 25410 38500
rect 11930 38420 25410 38430
rect 1890 30660 2000 35610
rect 4550 35010 4630 35610
rect 4530 35000 4650 35010
rect 4530 34930 4560 35000
rect 4620 34930 4650 35000
rect 4530 34920 4650 34930
rect 2070 33360 3000 33420
rect 2070 32670 2120 33360
rect 2950 32670 3000 33360
rect 2070 32620 3000 32670
rect 3100 33360 4030 33420
rect 3100 32670 3150 33360
rect 3980 32670 4030 33360
rect 3100 32620 4030 32670
rect 4130 33360 5060 33420
rect 4130 32670 4180 33360
rect 5010 32670 5060 33360
rect 4130 32620 5060 32670
rect 5160 33360 6090 33420
rect 5160 32670 5210 33360
rect 6040 32670 6090 33360
rect 5160 32620 6090 32670
rect 6190 33360 7120 33420
rect 6190 32670 6240 33360
rect 7070 32670 7120 33360
rect 6190 32620 7120 32670
rect 7220 33360 8150 33420
rect 7220 32670 7270 33360
rect 8100 32670 8150 33360
rect 7220 32620 8150 32670
rect 8250 33360 9180 33420
rect 8250 32670 8300 33360
rect 9130 32670 9180 33360
rect 8250 32620 9180 32670
rect 9280 33360 10920 33420
rect 9280 32670 9330 33360
rect 10870 32670 10920 33360
rect 9280 32620 10920 32670
rect 2070 32480 3000 32540
rect 2070 31790 2120 32480
rect 2950 31790 3000 32480
rect 2070 31740 3000 31790
rect 3100 32480 4030 32540
rect 3100 31790 3150 32480
rect 3980 31790 4030 32480
rect 3100 31740 4030 31790
rect 4130 32480 5060 32540
rect 4130 31790 4180 32480
rect 5010 31790 5060 32480
rect 4130 31740 5060 31790
rect 5160 32480 6090 32540
rect 5160 31790 5210 32480
rect 6040 31790 6090 32480
rect 5160 31740 6090 31790
rect 6190 32480 7120 32540
rect 6190 31790 6240 32480
rect 7070 31790 7120 32480
rect 6190 31740 7120 31790
rect 7220 32480 8150 32540
rect 7220 31790 7270 32480
rect 8100 31790 8150 32480
rect 7220 31740 8150 31790
rect 8250 32480 9180 32540
rect 8250 31790 8300 32480
rect 9130 31790 9180 32480
rect 8250 31740 9180 31790
rect 9280 32480 10210 32540
rect 9280 31790 9330 32480
rect 10160 31790 10210 32480
rect 9280 31740 10210 31790
rect 10310 32480 11240 32540
rect 10310 31790 10360 32480
rect 11190 31790 11240 32480
rect 10310 31740 11240 31790
rect 2930 30740 3050 30760
rect 2930 30680 2960 30740
rect 3020 30680 3050 30740
rect 2930 30670 3050 30680
rect 2930 30660 3040 30670
rect 1890 30580 3040 30660
rect 2070 29000 3000 29060
rect 2070 28310 2120 29000
rect 2950 28310 3000 29000
rect 2070 28260 3000 28310
rect 3100 29000 4030 29060
rect 3100 28310 3150 29000
rect 3980 28310 4030 29000
rect 3100 28260 4030 28310
rect 4130 29000 5060 29060
rect 4130 28310 4180 29000
rect 5010 28310 5060 29000
rect 4130 28260 5060 28310
rect 5160 29000 6090 29060
rect 5160 28310 5210 29000
rect 6040 28310 6090 29000
rect 5160 28260 6090 28310
rect 6190 29000 7120 29060
rect 6190 28310 6240 29000
rect 7070 28310 7120 29000
rect 6190 28260 7120 28310
rect 7220 29000 8150 29060
rect 7220 28310 7270 29000
rect 8100 28310 8150 29000
rect 7220 28260 8150 28310
rect 8250 29000 9180 29060
rect 8250 28310 8300 29000
rect 9130 28310 9180 29000
rect 8250 28260 9180 28310
rect 9280 29000 10210 29060
rect 9280 28310 9330 29000
rect 10160 28310 10210 29000
rect 9280 28260 10210 28310
rect 10310 29000 11240 29060
rect 10310 28310 10360 29000
rect 11190 28310 11240 29000
rect 10310 28260 11240 28310
rect 11930 28200 12020 38420
rect 25320 38410 25410 38420
rect 25620 37440 25700 44410
rect 25830 38510 25920 38520
rect 26170 38510 26250 44410
rect 25830 38500 26250 38510
rect 25830 38430 25840 38500
rect 25910 38430 26250 38500
rect 25830 38420 26250 38430
rect 25830 38410 25920 38420
rect 16350 37360 25700 37440
rect 12920 37200 13810 37260
rect 12920 36400 12970 37200
rect 13760 36400 13810 37200
rect 12920 36340 13810 36400
rect 13920 37200 14810 37260
rect 13920 36400 13970 37200
rect 14760 36400 14810 37200
rect 13920 36340 14810 36400
rect 16350 36160 16420 37360
rect 20710 36170 20810 36190
rect 20710 36160 20730 36170
rect 16350 36100 20730 36160
rect 15550 35630 15660 35640
rect 15550 35570 15570 35630
rect 15640 35620 15660 35630
rect 15760 35630 15930 35640
rect 15760 35620 15790 35630
rect 15640 35580 15790 35620
rect 15640 35570 15660 35580
rect 15550 35560 15660 35570
rect 15760 35570 15790 35580
rect 15900 35570 15930 35630
rect 15760 35560 15930 35570
rect 15790 34550 15900 35560
rect 16350 35510 16410 36100
rect 16350 35490 16530 35510
rect 16350 35430 16450 35490
rect 16510 35430 16530 35490
rect 16350 35410 16530 35430
rect 17220 35310 17330 35330
rect 17220 35240 17240 35310
rect 17310 35240 17330 35310
rect 17220 35220 17330 35240
rect 17970 34810 18020 36100
rect 20710 36090 20730 36100
rect 20790 36090 20810 36170
rect 20710 36070 20810 36090
rect 22230 36150 23290 36210
rect 22230 36040 22300 36150
rect 20410 35970 22300 36040
rect 18260 35300 18350 35320
rect 20410 35300 20480 35970
rect 20710 35910 20810 35930
rect 20710 35830 20730 35910
rect 20790 35830 20810 35910
rect 20710 35810 20810 35830
rect 18260 35230 18270 35300
rect 18340 35230 20480 35300
rect 18260 35210 18350 35230
rect 19730 34810 19830 34830
rect 17970 34750 19750 34810
rect 19810 34750 19830 34810
rect 19730 34730 19830 34750
rect 15420 34480 15900 34550
rect 18290 34620 18390 34630
rect 18290 34540 18310 34620
rect 18370 34540 18390 34620
rect 18290 34530 18390 34540
rect 14370 32010 14540 32020
rect 14370 31950 14400 32010
rect 14510 32000 14540 32010
rect 15420 32000 15480 34480
rect 19560 34430 19660 34450
rect 19560 34350 19580 34430
rect 19640 34350 19660 34430
rect 19560 34330 19660 34350
rect 15630 32310 15730 32340
rect 15630 32250 15650 32310
rect 15710 32250 15730 32310
rect 19580 32290 19640 34330
rect 20410 34320 20480 35230
rect 20730 34980 20790 35810
rect 22180 35310 22290 35330
rect 22180 35240 22200 35310
rect 22270 35240 22290 35310
rect 22180 35220 22290 35240
rect 23230 35280 23290 36150
rect 23230 35240 25510 35280
rect 23230 35230 23520 35240
rect 23510 35170 23520 35230
rect 23590 35230 25510 35240
rect 23590 35170 23600 35230
rect 23510 35150 23600 35170
rect 20730 34960 21000 34980
rect 20730 34900 20920 34960
rect 20980 34900 21000 34960
rect 20730 34880 21000 34900
rect 20740 34530 20840 34550
rect 20740 34450 20760 34530
rect 20820 34450 20840 34530
rect 20740 34430 20840 34450
rect 20410 34230 20720 34320
rect 15630 32220 15730 32250
rect 15930 32250 19640 32290
rect 15570 32020 15670 32040
rect 15570 32000 15590 32020
rect 14510 31960 15590 32000
rect 14510 31950 14540 31960
rect 14370 31940 14540 31950
rect 15570 31940 15590 31960
rect 15650 31940 15670 32020
rect 15570 31920 15670 31940
rect 15930 31470 15970 32250
rect 15930 31450 16530 31470
rect 15930 31390 16450 31450
rect 16510 31390 16530 31450
rect 15930 31370 16530 31390
rect 17220 31300 17330 31320
rect 17220 31230 17240 31300
rect 17310 31230 17330 31300
rect 17220 31210 17330 31230
rect 20640 31170 20720 34230
rect 18530 31150 20720 31170
rect 18530 31080 18540 31150
rect 18610 31100 20720 31150
rect 18610 31080 18620 31100
rect 18530 31060 18620 31080
rect 20750 30860 20820 34430
rect 20900 34410 21000 34880
rect 24690 34810 24790 34830
rect 24620 34750 24710 34810
rect 24770 34750 24790 34810
rect 23220 34550 23320 34560
rect 23220 34470 23240 34550
rect 23300 34470 23320 34550
rect 23220 34460 23320 34470
rect 20900 34370 22380 34410
rect 20900 34320 21000 34370
rect 20720 30840 20820 30860
rect 19990 30750 20090 30770
rect 19990 30690 20010 30750
rect 20070 30690 20090 30750
rect 20720 30760 20740 30840
rect 20800 30760 20820 30840
rect 20720 30740 20820 30760
rect 20870 34250 21000 34320
rect 22340 34280 22380 34370
rect 22740 34380 24220 34420
rect 22740 34280 22780 34380
rect 19990 30660 20090 30690
rect 20870 30660 20920 34250
rect 22340 34240 22780 34280
rect 24180 34300 24220 34380
rect 24620 34300 24660 34750
rect 24690 34730 24790 34750
rect 24180 34260 24660 34300
rect 24930 34380 25030 34400
rect 24930 34300 24950 34380
rect 25010 34300 25030 34380
rect 24930 34280 25030 34300
rect 22390 34060 23130 34120
rect 22390 33250 22440 34060
rect 23080 33250 23130 34060
rect 24950 34040 25010 34280
rect 22390 33190 23130 33250
rect 24450 33980 25010 34040
rect 24450 32360 24510 33980
rect 20990 32320 24510 32360
rect 20990 30920 21040 32320
rect 25440 31390 25510 35230
rect 25180 31330 25510 31390
rect 22240 31300 22350 31320
rect 22240 31230 22260 31300
rect 22330 31230 22350 31300
rect 22240 31210 22350 31230
rect 25180 31170 25250 31330
rect 23560 31150 25250 31170
rect 23560 31080 23570 31150
rect 23640 31100 25250 31150
rect 23640 31080 23650 31100
rect 23560 31060 23650 31080
rect 20960 30900 21060 30920
rect 20960 30840 20980 30900
rect 21040 30840 21060 30900
rect 20960 30820 21060 30840
rect 24950 30740 25050 30760
rect 19990 30620 20920 30660
rect 18220 30480 18330 30490
rect 18220 30400 18240 30480
rect 18310 30400 18330 30480
rect 18220 30390 18330 30400
rect 20540 30460 20640 30480
rect 20540 30380 20560 30460
rect 20620 30380 20640 30460
rect 15380 30280 15490 30300
rect 15380 30210 15400 30280
rect 15470 30210 15490 30280
rect 15380 30190 15490 30210
rect 12700 28620 12840 28640
rect 12700 28510 12720 28620
rect 12820 28510 12840 28620
rect 12700 28490 12840 28510
rect 6280 28130 12020 28200
rect 12690 28270 12830 28290
rect 12690 28160 12710 28270
rect 12810 28160 12830 28270
rect 12690 28140 12830 28160
rect 5360 28100 5500 28120
rect 5360 27990 5380 28100
rect 5480 27990 5500 28100
rect 5360 27970 5500 27990
rect 5590 27820 5730 27840
rect 5590 27710 5610 27820
rect 5710 27710 5730 27820
rect 5590 27690 5730 27710
rect 6280 25560 6380 28130
rect 20540 27690 20640 30380
rect 6280 25500 6300 25560
rect 6360 25500 6380 25560
rect 6280 25480 6380 25500
rect 6430 27610 20640 27690
rect 20720 30460 20820 30480
rect 20720 30380 20740 30460
rect 20800 30380 20820 30460
rect 6430 18700 6510 27610
rect 20720 27570 20820 30380
rect 20870 30340 20920 30620
rect 24880 30680 24970 30740
rect 25030 30680 25050 30740
rect 23240 30480 23340 30490
rect 23240 30400 23260 30480
rect 23320 30400 23340 30480
rect 23240 30390 23340 30400
rect 20870 30300 22440 30340
rect 22400 30210 22440 30300
rect 22800 30310 24280 30350
rect 22800 30210 22840 30310
rect 22400 30170 22840 30210
rect 24240 30230 24280 30310
rect 24880 30230 24920 30680
rect 24950 30660 25050 30680
rect 24240 30190 24920 30230
rect 22390 29980 23130 30040
rect 22390 29170 22440 29980
rect 23080 29170 23130 29980
rect 22390 29110 23130 29170
rect 6560 27480 20820 27570
rect 6560 19490 6640 27480
rect 7320 27360 8250 27420
rect 7320 26670 7370 27360
rect 8200 26670 8250 27360
rect 7320 26620 8250 26670
rect 8350 27360 9280 27420
rect 8350 26670 8400 27360
rect 9230 26670 9280 27360
rect 8350 26620 9280 26670
rect 9380 27360 10310 27420
rect 9380 26670 9430 27360
rect 10260 26670 10310 27360
rect 9380 26620 10310 26670
rect 10410 27360 11340 27420
rect 10410 26670 10460 27360
rect 11290 26670 11340 27360
rect 10410 26620 11340 26670
rect 11440 27360 12370 27420
rect 11440 26670 11490 27360
rect 12320 26670 12370 27360
rect 11440 26620 12370 26670
rect 12470 27360 13400 27420
rect 12470 26670 12520 27360
rect 13350 26670 13400 27360
rect 12470 26620 13400 26670
rect 13500 27360 14430 27420
rect 13500 26670 13550 27360
rect 14380 26670 14430 27360
rect 13500 26620 14430 26670
rect 14530 27360 15460 27420
rect 14530 26670 14580 27360
rect 15410 26670 15460 27360
rect 14530 26620 15460 26670
rect 15560 27360 16490 27420
rect 15560 26670 15610 27360
rect 16440 26670 16490 27360
rect 15560 26620 16490 26670
rect 16590 27360 17520 27420
rect 16590 26670 16640 27360
rect 17470 26670 17520 27360
rect 16590 26620 17520 26670
rect 17620 27360 18550 27420
rect 17620 26670 17670 27360
rect 18500 26670 18550 27360
rect 17620 26620 18550 26670
rect 18650 27360 19580 27420
rect 18650 26670 18700 27360
rect 19530 26670 19580 27360
rect 18650 26620 19580 26670
rect 19710 27360 20640 27420
rect 19710 26670 19760 27360
rect 20590 26670 20640 27360
rect 19710 26620 20640 26670
rect 8350 26460 11480 26520
rect 7420 24870 8160 24880
rect 7420 24820 8080 24870
rect 6560 19470 7190 19490
rect 6560 19410 7110 19470
rect 7170 19410 7190 19470
rect 6560 19390 7190 19410
rect 6430 18680 7290 18700
rect 6430 18620 6960 18680
rect 7020 18620 7290 18680
rect 6430 18600 7290 18620
rect 7230 18440 7290 18600
rect 7210 18420 7310 18440
rect 7210 18360 7230 18420
rect 7290 18360 7310 18420
rect 7210 18340 7310 18360
rect 7420 15310 7500 24820
rect 8060 24800 8080 24820
rect 8140 24800 8160 24870
rect 8060 24790 8160 24800
rect 7530 24770 7650 24790
rect 7530 24710 7570 24770
rect 7630 24730 7760 24770
rect 8180 24730 8280 24750
rect 7630 24710 8200 24730
rect 7530 24690 7650 24710
rect 7700 24670 8200 24710
rect 8260 24670 8280 24730
rect 7700 22790 7760 24670
rect 8180 24650 8280 24670
rect 8350 23140 8410 26460
rect 11410 24870 11480 26460
rect 10400 24850 10490 24870
rect 10400 24790 10410 24850
rect 10480 24790 10490 24850
rect 10400 24770 10490 24790
rect 11400 24850 11490 24870
rect 11400 24790 11410 24850
rect 11480 24790 11490 24850
rect 11400 24770 11490 24790
rect 10410 24700 10480 24770
rect 10410 24640 10520 24700
rect 9080 24440 9170 24460
rect 9080 24380 9090 24440
rect 9160 24380 9170 24440
rect 9080 24360 9170 24380
rect 9090 24140 9160 24360
rect 10470 24140 10520 24640
rect 9090 24060 10520 24140
rect 9080 23140 9170 23160
rect 8350 23080 9090 23140
rect 9160 23080 9170 23140
rect 9080 23060 9170 23080
rect 10470 22910 10520 24060
rect 19500 24190 20430 24240
rect 19500 23380 19560 24190
rect 20370 23380 20430 24190
rect 19500 23330 20430 23380
rect 10410 22870 10520 22910
rect 10410 22800 10480 22870
rect 7700 22730 9290 22790
rect 9100 18330 9170 22730
rect 9200 22700 9290 22730
rect 10400 22780 10490 22800
rect 10400 22720 10410 22780
rect 10480 22720 10490 22780
rect 10400 22700 10490 22720
rect 11400 22780 11490 22800
rect 11400 22720 11410 22780
rect 11480 22720 11490 22780
rect 11400 22700 11490 22720
rect 9200 22640 9220 22700
rect 9280 22640 9290 22700
rect 9200 22620 9290 22640
rect 9200 18330 9290 18350
rect 9100 18270 9220 18330
rect 9280 18270 9290 18330
rect 10410 18280 10480 22700
rect 9200 18250 9290 18270
rect 10400 18260 10490 18280
rect 10400 18200 10410 18260
rect 10480 18200 10490 18260
rect 10400 18180 10490 18200
rect 9460 18100 9550 18120
rect 8430 18040 9470 18100
rect 9540 18040 9550 18100
rect 7420 15290 7510 15310
rect 7420 15230 7430 15290
rect 7500 15230 7510 15290
rect 7420 15210 7510 15230
rect 7420 13000 7500 15210
rect 8430 14280 8500 18040
rect 9460 18020 9550 18040
rect 9080 17960 9170 17980
rect 9080 17900 9090 17960
rect 9160 17900 9170 17960
rect 9080 17880 9170 17900
rect 9090 17840 9140 17880
rect 11430 17840 11480 22700
rect 17620 20890 18550 20950
rect 12720 20410 12810 20430
rect 12720 20350 12730 20410
rect 12800 20350 13020 20410
rect 12720 20330 12810 20350
rect 9090 17790 11480 17840
rect 12950 16700 13020 20350
rect 17620 20090 17670 20890
rect 18500 20090 18550 20890
rect 17620 20030 18550 20090
rect 19500 17600 20430 17650
rect 19500 16790 19560 17600
rect 20370 16790 20430 17600
rect 19500 16740 20430 16790
rect 10660 16630 13020 16700
rect 10660 15810 10730 16630
rect 10170 15740 10730 15810
rect 10870 16410 11800 16470
rect 9670 15110 9830 15120
rect 9670 15050 9750 15110
rect 9810 15050 9830 15110
rect 9670 15040 9830 15050
rect 8420 14260 8510 14280
rect 8420 14200 8430 14260
rect 8500 14200 8510 14260
rect 8420 14180 8510 14200
rect 9670 13170 9720 15040
rect 10170 15030 10240 15740
rect 10870 15720 10920 16410
rect 11750 15720 11800 16410
rect 10870 15670 11800 15720
rect 11900 16410 12830 16470
rect 11900 15720 11950 16410
rect 12780 15720 12830 16410
rect 11900 15670 12830 15720
rect 12930 16410 13860 16470
rect 12930 15720 12980 16410
rect 13810 15720 13860 16410
rect 12930 15670 13860 15720
rect 13990 16410 14920 16470
rect 13990 15720 14040 16410
rect 14870 15720 14920 16410
rect 13990 15670 14920 15720
rect 15020 16410 15950 16470
rect 15020 15720 15070 16410
rect 15900 15720 15950 16410
rect 15020 15670 15950 15720
rect 16050 16410 16980 16470
rect 16050 15720 16100 16410
rect 16930 15720 16980 16410
rect 16050 15670 16980 15720
rect 17110 16410 18040 16470
rect 17110 15720 17160 16410
rect 17990 15720 18040 16410
rect 17110 15670 18040 15720
rect 18140 16410 19070 16470
rect 18140 15720 18190 16410
rect 19020 15720 19070 16410
rect 18140 15670 19070 15720
rect 19170 16410 20100 16470
rect 19170 15720 19220 16410
rect 20050 15720 20100 16410
rect 19170 15670 20100 15720
rect 20230 16410 21160 16470
rect 20230 15720 20280 16410
rect 21110 15720 21160 16410
rect 20230 15670 21160 15720
rect 10170 15020 10370 15030
rect 10170 14960 10280 15020
rect 10350 14960 10370 15020
rect 10170 14950 10370 14960
rect 9850 14240 10780 14290
rect 9850 13430 9910 14240
rect 10720 13430 10780 14240
rect 9850 13380 10780 13430
rect 10880 14240 11810 14290
rect 10880 13430 10940 14240
rect 11750 13430 11810 14240
rect 10880 13380 11810 13430
rect 11910 14240 12840 14290
rect 11910 13430 11970 14240
rect 12780 13430 12840 14240
rect 11910 13380 12840 13430
rect 12920 14240 13850 14290
rect 12920 13430 12980 14240
rect 13790 13430 13850 14240
rect 12920 13380 13850 13430
rect 9660 13150 9750 13170
rect 9660 13090 9670 13150
rect 9740 13090 9750 13150
rect 9660 13070 9750 13090
rect 7420 12930 11350 13000
rect 7640 12710 7800 12720
rect 7640 12650 7700 12710
rect 7760 12650 7800 12710
rect 7640 12640 7800 12650
rect 7570 12600 7670 12610
rect 7570 12540 7590 12600
rect 7650 12540 7670 12600
rect 7570 12530 7670 12540
rect 7600 10960 7650 12530
rect 7590 10950 7690 10960
rect 7590 10890 7610 10950
rect 7670 10890 7690 10950
rect 7590 10880 7690 10890
rect 7720 10850 7780 12640
rect 11290 12630 11350 12930
rect 11270 12610 11360 12630
rect 11270 12550 11280 12610
rect 11350 12550 11360 12610
rect 9740 12530 9830 12550
rect 11270 12530 11360 12550
rect 9740 12470 9750 12530
rect 9820 12470 9830 12530
rect 9740 12450 9830 12470
rect 9770 10950 9830 12450
rect 9650 10900 9830 10950
rect 7840 10850 7920 10870
rect 9650 10860 9720 10900
rect 7720 10790 7850 10850
rect 7910 10790 7920 10850
rect 7840 10770 7920 10790
rect 9630 10840 9740 10860
rect 9630 10780 9650 10840
rect 9720 10780 9740 10840
rect 9630 10760 9740 10780
rect 11290 10550 11340 12530
rect 13990 11860 14920 11920
rect 13990 11170 14040 11860
rect 14870 11170 14920 11860
rect 13990 11120 14920 11170
rect 15020 11860 15950 11920
rect 15020 11170 15070 11860
rect 15900 11170 15950 11860
rect 15020 11120 15950 11170
rect 16050 11860 16980 11920
rect 16050 11170 16100 11860
rect 16930 11170 16980 11860
rect 16050 11120 16980 11170
rect 17110 11860 18040 11920
rect 17110 11170 17160 11860
rect 17990 11170 18040 11860
rect 17110 11120 18040 11170
rect 18140 11860 19070 11920
rect 18140 11170 18190 11860
rect 19020 11170 19070 11860
rect 18140 11120 19070 11170
rect 19170 11860 20100 11920
rect 19170 11170 19220 11860
rect 20050 11170 20100 11860
rect 19170 11120 20100 11170
rect 20230 11860 21160 11920
rect 20230 11170 20280 11860
rect 21110 11170 21160 11860
rect 20230 11120 21160 11170
rect 11280 10530 11370 10550
rect 11280 10470 11290 10530
rect 11360 10470 11370 10530
rect 11280 10450 11370 10470
rect 12280 10500 12370 10520
rect 12280 10440 12290 10500
rect 12360 10440 12370 10500
rect 9770 10410 9880 10430
rect 12280 10420 12370 10440
rect 9770 10350 9790 10410
rect 9860 10350 9880 10410
rect 9770 10330 9880 10350
rect 9800 9780 9850 10330
rect 12290 9780 12360 10420
rect 9800 9740 12360 9780
rect 8820 9610 9750 9670
rect 8820 8800 8880 9610
rect 9690 8800 9750 9610
rect 8820 8750 9750 8800
rect 9850 9610 10780 9670
rect 9850 8800 9910 9610
rect 10720 8800 10780 9610
rect 9850 8750 10780 8800
rect 10880 9610 11810 9670
rect 10880 8800 10940 9610
rect 11750 8800 11810 9610
rect 10880 8750 11810 8800
rect 11910 9610 12840 9670
rect 11910 8800 11970 9610
rect 12780 8800 12840 9610
rect 11910 8750 12840 8800
rect 12920 9610 13850 9670
rect 12920 8800 12980 9610
rect 13790 8800 13850 9610
rect 12920 8750 13850 8800
rect 13950 9610 14880 9670
rect 13950 8800 14010 9610
rect 14820 8800 14880 9610
rect 13950 8750 14880 8800
rect 14980 9610 15910 9670
rect 14980 8800 15040 9610
rect 15850 8800 15910 9610
rect 14980 8750 15910 8800
rect 16010 9610 16940 9670
rect 16010 8800 16070 9610
rect 16880 8800 16940 9610
rect 16010 8750 16940 8800
rect 17020 9610 17950 9670
rect 17020 8800 17080 9610
rect 17890 8800 17950 9610
rect 17020 8750 17950 8800
rect 18050 9610 18980 9670
rect 18050 8800 18110 9610
rect 18920 8800 18980 9610
rect 18050 8750 18980 8800
rect 19060 9610 19990 9670
rect 19060 8800 19120 9610
rect 19930 8800 19990 9610
rect 19060 8750 19990 8800
rect 20090 9610 21160 9670
rect 20090 8800 20150 9610
rect 21110 8800 21160 9610
rect 21550 8920 21660 8940
rect 21550 8850 21570 8920
rect 21640 8850 21660 8920
rect 21550 8830 21660 8850
rect 21950 8920 22060 8940
rect 21950 8850 21970 8920
rect 22040 8850 22060 8920
rect 21950 8830 22060 8850
rect 22380 8920 22490 8940
rect 22380 8850 22400 8920
rect 22470 8850 22490 8920
rect 22380 8830 22490 8850
rect 20090 8750 21160 8800
rect 13390 8490 13600 8510
rect 13390 8420 13430 8490
rect 13560 8420 13600 8490
rect 13390 8400 13600 8420
rect 9870 6870 11260 6920
rect 9870 6060 9930 6870
rect 11200 6060 11260 6870
rect 9870 6000 11260 6060
rect 11370 6870 12300 6920
rect 11370 6060 11430 6870
rect 12240 6060 12300 6870
rect 11370 6000 12300 6060
rect 12400 6870 13330 6920
rect 12400 6060 12460 6870
rect 13270 6060 13330 6870
rect 12400 6000 13330 6060
rect 13430 5900 13510 8400
rect 13600 6870 14990 6920
rect 13600 6060 13660 6870
rect 14930 6060 14990 6870
rect 13600 6000 14990 6060
rect 15100 6870 16030 6920
rect 15100 6060 15160 6870
rect 15970 6060 16030 6870
rect 15100 6000 16030 6060
rect 16130 6870 17060 6920
rect 16130 6060 16190 6870
rect 17000 6060 17060 6870
rect 16130 6000 17060 6060
rect 13340 5880 13550 5900
rect 13340 5820 13380 5880
rect 13510 5820 13550 5880
rect 13340 5800 13550 5820
rect 13340 4500 13550 4520
rect 13340 4440 13380 4500
rect 13510 4440 13550 4500
rect 13340 4420 13550 4440
rect 13340 4340 13550 4360
rect 13340 4280 13380 4340
rect 13510 4280 13550 4340
rect 13340 4260 13550 4280
rect 19180 4170 19330 4200
rect 9840 4140 9940 4160
rect 9840 4070 9850 4140
rect 9930 4070 9940 4140
rect 9840 4050 9940 4070
rect 19180 4070 19200 4170
rect 19310 4070 19330 4170
rect 19180 4040 19330 4070
rect 200 3990 600 4010
rect 200 3880 230 3990
rect 570 3880 600 3990
rect 200 3860 600 3880
rect 13280 3080 13490 3100
rect 13280 3020 13320 3080
rect 13450 3020 13490 3080
rect 13280 3000 13490 3020
rect 9850 2840 11190 2890
rect 9850 2030 9910 2840
rect 11130 2030 11190 2840
rect 9850 1980 11190 2030
rect 11290 2840 12220 2890
rect 11290 2030 11350 2840
rect 12160 2030 12220 2840
rect 11290 1980 12220 2030
rect 12310 2840 13240 2890
rect 12310 2030 12370 2840
rect 13180 2030 13240 2840
rect 12310 1980 13240 2030
rect 13350 620 13450 3000
rect 13510 2840 15010 2890
rect 13510 2030 13570 2840
rect 14950 2030 15010 2840
rect 13510 1980 15010 2030
rect 15110 2840 16040 2890
rect 15110 2030 15170 2840
rect 15980 2030 16040 2840
rect 15110 1980 16040 2030
rect 16130 2840 17060 2890
rect 16130 2030 16190 2840
rect 17000 2030 17060 2840
rect 16130 1980 17060 2030
rect 13320 600 13530 620
rect 13320 530 13360 600
rect 13490 530 13530 600
rect 13320 510 13530 530
rect 21570 440 21640 8830
rect 21970 4330 22040 8830
rect 22400 4330 22470 8830
rect 22550 8640 22660 8660
rect 23250 8640 23360 8660
rect 22550 8570 22570 8640
rect 22640 8570 23270 8640
rect 23340 8570 23360 8640
rect 22550 8550 22660 8570
rect 23250 8550 23360 8570
rect 21950 4310 22060 4330
rect 21950 4240 21970 4310
rect 22040 4240 22060 4310
rect 21950 4220 22060 4240
rect 22380 4310 22490 4330
rect 22380 4240 22400 4310
rect 22470 4240 22490 4310
rect 22380 4220 22490 4240
rect 27200 2780 27600 2810
rect 23110 2710 24210 2770
rect 23110 2080 23170 2710
rect 23980 2080 24210 2710
rect 27200 2130 27230 2780
rect 27570 2130 27600 2780
rect 27200 2100 27600 2130
rect 23110 2030 24210 2080
rect 21550 420 21660 440
rect 21550 350 21570 420
rect 21640 350 21660 420
rect 21550 330 21660 350
<< via2 >>
rect 24520 44430 24600 44560
rect 2120 43410 2950 44100
rect 3430 42310 4280 43000
rect 10060 39880 10900 40000
rect 2130 38620 3170 39430
rect 3380 38620 4420 39430
rect 4630 38620 5670 39430
rect 5880 38620 6920 39430
rect 7130 38620 8170 39430
rect 8380 38620 9850 39430
rect 2120 37240 3860 38050
rect 4070 37240 5110 38050
rect 5320 37240 6360 38050
rect 6570 37240 7610 38050
rect 7820 37240 8860 38050
rect 9070 37240 9820 38050
rect 10080 37240 10880 38050
rect 25620 44430 25700 44560
rect 26170 44430 26250 44560
rect 21730 43410 22580 44100
rect 22980 43410 23830 44100
rect 15690 43050 15770 43180
rect 23640 41810 23720 41870
rect 21610 40340 22250 41020
rect 22440 40340 23080 41020
rect 23260 40340 23900 41020
rect 2120 32670 2950 33360
rect 3150 32670 3980 33360
rect 4180 32670 5010 33360
rect 5210 32670 6040 33360
rect 6240 32670 7070 33360
rect 7270 32670 8100 33360
rect 8300 32670 9130 33360
rect 9330 32670 10870 33360
rect 2120 31790 2950 32480
rect 3150 31790 3980 32480
rect 4180 31790 5010 32480
rect 5210 31790 6040 32480
rect 6240 31790 7070 32480
rect 7270 31790 8100 32480
rect 8300 31790 9130 32480
rect 9330 31790 10160 32480
rect 10360 31790 11190 32480
rect 2120 28310 2950 29000
rect 3150 28310 3980 29000
rect 4180 28310 5010 29000
rect 5210 28310 6040 29000
rect 6240 28310 7070 29000
rect 7270 28310 8100 29000
rect 8300 28310 9130 29000
rect 9330 28310 10160 29000
rect 10360 28310 11190 29000
rect 12970 36400 13760 37200
rect 13970 36400 14760 37200
rect 17240 35240 17310 35310
rect 18310 34540 18370 34620
rect 15650 32250 15710 32310
rect 22200 35240 22270 35310
rect 17240 31230 17310 31300
rect 23240 34470 23300 34550
rect 22440 33250 23080 34060
rect 22260 31230 22330 31300
rect 18240 30400 18310 30480
rect 15400 30210 15470 30280
rect 12720 28510 12820 28620
rect 12710 28160 12810 28270
rect 5380 27990 5480 28100
rect 5610 27710 5710 27820
rect 23260 30400 23320 30480
rect 22440 29170 23080 29980
rect 7370 26670 8200 27360
rect 8400 26670 9230 27360
rect 9430 26670 10260 27360
rect 10460 26670 11290 27360
rect 11490 26670 12320 27360
rect 12520 26670 13350 27360
rect 13550 26670 14380 27360
rect 14580 26670 15410 27360
rect 15610 26670 16440 27360
rect 16640 26670 17470 27360
rect 17670 26670 18500 27360
rect 18700 26670 19530 27360
rect 19760 26670 20590 27360
rect 19560 23380 20370 24190
rect 17670 20090 18500 20890
rect 19560 16790 20370 17600
rect 10920 15720 11750 16410
rect 11950 15720 12780 16410
rect 12980 15720 13810 16410
rect 14040 15720 14870 16410
rect 15070 15720 15900 16410
rect 16100 15720 16930 16410
rect 17160 15720 17990 16410
rect 18190 15720 19020 16410
rect 19220 15720 20050 16410
rect 20280 15720 21110 16410
rect 9910 13430 10720 14240
rect 10940 13430 11750 14240
rect 11970 13430 12780 14240
rect 12980 13430 13790 14240
rect 14040 11170 14870 11860
rect 15070 11170 15900 11860
rect 16100 11170 16930 11860
rect 17160 11170 17990 11860
rect 18190 11170 19020 11860
rect 19220 11170 20050 11860
rect 20280 11170 21110 11860
rect 8880 8800 9690 9610
rect 9910 8800 10720 9610
rect 10940 8800 11750 9610
rect 11970 8800 12780 9610
rect 12980 8800 13790 9610
rect 14010 8800 14820 9610
rect 15040 8800 15850 9610
rect 16070 8800 16880 9610
rect 17080 8800 17890 9610
rect 18110 8800 18920 9610
rect 19120 8800 19930 9610
rect 20150 8800 21110 9610
rect 9930 6060 11200 6870
rect 11430 6060 12240 6870
rect 12460 6060 13270 6870
rect 13660 6060 14930 6870
rect 15160 6060 15970 6870
rect 16190 6060 17000 6870
rect 9850 4070 9930 4140
rect 19200 4070 19310 4170
rect 230 3880 570 3990
rect 9910 2030 11130 2840
rect 11350 2030 12160 2840
rect 12370 2030 13180 2840
rect 13570 2030 14950 2840
rect 15170 2030 15980 2840
rect 16190 2030 17000 2840
rect 23170 2080 23980 2710
rect 27230 2130 27570 2780
<< metal3 >>
rect 24500 44560 24620 44580
rect 24500 44430 24520 44560
rect 24600 44430 24620 44560
rect 24500 44410 24620 44430
rect 25600 44560 25720 44580
rect 25600 44430 25620 44560
rect 25700 44430 25720 44560
rect 25600 44410 25720 44430
rect 26150 44560 26270 44580
rect 26150 44430 26170 44560
rect 26250 44430 26270 44560
rect 26150 44410 26270 44430
rect 200 44130 23880 44160
rect 200 44120 12950 44130
rect 200 43390 230 44120
rect 570 44100 12950 44120
rect 570 43410 2120 44100
rect 2950 43410 12950 44100
rect 570 43390 12950 43410
rect 13780 44120 23880 44130
rect 13780 43390 13950 44120
rect 200 43380 13950 43390
rect 14780 44100 23880 44120
rect 14780 43410 21730 44100
rect 22580 43410 22980 44100
rect 23830 43410 23880 44100
rect 14780 43380 23880 43410
rect 200 43360 23880 43380
rect 15670 43180 15790 43200
rect 800 43030 4330 43060
rect 15670 43050 15690 43180
rect 15770 43050 15790 43180
rect 15670 43030 15790 43050
rect 800 42290 830 43030
rect 1170 43000 4330 43030
rect 1170 42310 3430 43000
rect 4280 42310 4330 43000
rect 1170 42290 4330 42310
rect 800 42260 4330 42290
rect 11720 41880 23740 41890
rect 11720 41800 11740 41880
rect 11820 41870 23740 41880
rect 11820 41810 23640 41870
rect 23720 41810 23740 41870
rect 11820 41800 23740 41810
rect 11720 41790 23740 41800
rect 800 41050 23950 41080
rect 800 40320 830 41050
rect 1170 41020 23950 41050
rect 1170 40340 21610 41020
rect 22250 40340 22440 41020
rect 23080 40340 23260 41020
rect 23900 40340 23950 41020
rect 1170 40320 23950 40340
rect 800 40290 23950 40320
rect 10030 40000 10930 40020
rect 10030 39880 10060 40000
rect 10900 39880 10930 40000
rect 10030 39860 10930 39880
rect 10030 39830 27600 39860
rect 800 39460 9900 39490
rect 800 38590 830 39460
rect 1170 39430 9900 39460
rect 1170 38620 2130 39430
rect 3170 38620 3380 39430
rect 4420 38620 4630 39430
rect 5670 38620 5880 39430
rect 6920 38620 7130 39430
rect 8170 38620 8380 39430
rect 9850 38620 9900 39430
rect 10030 38900 10060 39830
rect 10900 38900 27230 39830
rect 27570 38900 27600 39830
rect 10030 38870 27600 38900
rect 1170 38590 9900 38620
rect 800 38560 9900 38590
rect 2070 38050 10930 38110
rect 2070 37240 2120 38050
rect 3860 37240 4070 38050
rect 5110 37240 5320 38050
rect 6360 37240 6570 38050
rect 7610 37240 7820 38050
rect 8860 37240 9070 38050
rect 9820 37240 10080 38050
rect 10880 37240 10930 38050
rect 2070 37180 10930 37240
rect 12920 37200 13810 37260
rect 12920 36400 12970 37200
rect 13760 36400 13810 37200
rect 12920 36340 13810 36400
rect 13920 37200 14810 37260
rect 13920 36400 13970 37200
rect 14760 36400 14810 37200
rect 13920 36340 14810 36400
rect 13880 34970 14940 35530
rect 17220 35310 17330 35330
rect 17220 35240 17240 35310
rect 17310 35240 17330 35310
rect 17220 35220 17330 35240
rect 20170 34970 21230 35650
rect 22180 35310 22290 35330
rect 22180 35240 22200 35310
rect 22270 35240 22290 35310
rect 22180 35220 22290 35240
rect 13880 34690 21370 34970
rect 13880 34500 15350 34690
rect 13880 34470 14940 34500
rect 1400 33390 10920 33420
rect 1400 32650 1430 33390
rect 1770 33360 10920 33390
rect 1770 32670 2120 33360
rect 2950 32670 3150 33360
rect 3980 32670 4180 33360
rect 5010 32670 5210 33360
rect 6040 32670 6240 33360
rect 7070 32670 7270 33360
rect 8100 32670 8300 33360
rect 9130 32670 9330 33360
rect 10870 32670 10920 33360
rect 1770 32650 10920 32670
rect 1400 32620 10920 32650
rect 800 32510 11240 32540
rect 800 31770 830 32510
rect 1170 32480 11240 32510
rect 1170 31790 2120 32480
rect 2950 31790 3150 32480
rect 3980 31790 4180 32480
rect 5010 31790 5210 32480
rect 6040 31790 6240 32480
rect 7070 31790 7270 32480
rect 8100 31790 8300 32480
rect 9130 31790 9330 32480
rect 10160 31790 10360 32480
rect 11190 31790 11240 32480
rect 1170 31770 11240 31790
rect 800 31740 11240 31770
rect 15100 31300 15350 34500
rect 18290 34620 18390 34630
rect 18290 34540 18310 34620
rect 18370 34540 18390 34620
rect 20170 34620 21370 34690
rect 20170 34590 21230 34620
rect 18290 34330 18390 34540
rect 23220 34550 23320 34560
rect 23220 34470 23240 34550
rect 23300 34470 23320 34550
rect 23220 34330 23320 34470
rect 15630 34250 23340 34330
rect 15630 32310 15730 34250
rect 22390 34060 23130 34120
rect 22390 33250 22440 34060
rect 23080 33250 23130 34060
rect 22390 33190 23130 33250
rect 15630 32250 15650 32310
rect 15710 32250 15730 32310
rect 15630 32220 15730 32250
rect 13620 30540 14680 31210
rect 15090 30850 15350 31300
rect 17220 31300 17330 31320
rect 17220 31230 17240 31300
rect 17310 31230 17330 31300
rect 17220 31210 17330 31230
rect 20180 31300 21240 31970
rect 22240 31300 22350 31320
rect 20180 30850 21660 31300
rect 22240 31230 22260 31300
rect 22330 31230 22350 31300
rect 22240 31210 22350 31230
rect 15100 30650 15350 30850
rect 21320 30650 21660 30850
rect 15100 30580 21660 30650
rect 15100 30540 15490 30580
rect 13620 30280 15490 30540
rect 23240 30490 23340 34250
rect 18220 30480 23340 30490
rect 18220 30400 18240 30480
rect 18310 30400 23260 30480
rect 23320 30400 23340 30480
rect 18220 30390 23340 30400
rect 13620 30230 15400 30280
rect 13620 30150 14680 30230
rect 15380 30210 15400 30230
rect 15470 30210 15490 30280
rect 15380 30190 15490 30210
rect 22390 29980 23130 30040
rect 22390 29170 22440 29980
rect 23080 29170 23130 29980
rect 22390 29110 23130 29170
rect 200 29030 11240 29060
rect 200 28290 230 29030
rect 570 29000 11240 29030
rect 570 28310 2120 29000
rect 2950 28310 3150 29000
rect 3980 28310 4180 29000
rect 5010 28310 5210 29000
rect 6040 28310 6240 29000
rect 7070 28310 7270 29000
rect 8100 28310 8300 29000
rect 9130 28310 9330 29000
rect 10160 28310 10360 29000
rect 11190 28310 11240 29000
rect 570 28290 11240 28310
rect 200 28260 11240 28290
rect 12260 28620 12840 28640
rect 12260 28510 12720 28620
rect 12820 28510 12840 28620
rect 12260 28490 12840 28510
rect 5360 28100 5500 28120
rect 12260 28100 12380 28490
rect 5360 27990 5380 28100
rect 5480 27990 12380 28100
rect 12690 28270 12830 28290
rect 12690 28160 12710 28270
rect 12810 28160 12830 28270
rect 5360 27970 5500 27990
rect 5590 27820 5730 27840
rect 12690 27820 12830 28160
rect 5590 27710 5610 27820
rect 5710 27710 12830 27820
rect 5590 27690 5730 27710
rect 1400 27400 20640 27430
rect 1400 26630 1430 27400
rect 1770 27360 20640 27400
rect 1770 26670 7370 27360
rect 8200 26670 8400 27360
rect 9230 26670 9430 27360
rect 10260 26670 10460 27360
rect 11290 26670 11490 27360
rect 12320 26670 12520 27360
rect 13350 26670 13550 27360
rect 14380 26670 14580 27360
rect 15410 26670 15610 27360
rect 16440 26910 16640 27360
rect 16440 26670 16490 26910
rect 1770 26630 16490 26670
rect 1400 26620 16490 26630
rect 16590 26670 16640 26910
rect 17470 26670 17670 27360
rect 18500 26670 18700 27360
rect 19530 26670 19760 27360
rect 20590 26670 20640 27360
rect 16590 26620 20640 26670
rect 1400 26600 15910 26620
rect 17020 26600 20640 26620
rect 17620 20890 18550 26600
rect 17620 20090 17670 20890
rect 18500 20090 18550 20890
rect 17620 20030 18550 20090
rect 19500 24210 27600 24240
rect 19500 24190 27230 24210
rect 19500 23380 19560 24190
rect 20370 23380 27230 24190
rect 19500 23360 27230 23380
rect 27570 23360 27600 24210
rect 19500 23330 27600 23360
rect 19500 17600 20430 23330
rect 19500 16790 19560 17600
rect 20370 16790 20430 17600
rect 19500 16740 20430 16790
rect 800 16440 21160 16470
rect 800 15700 830 16440
rect 1170 16410 21160 16440
rect 1170 15720 10920 16410
rect 11750 15720 11950 16410
rect 12780 15720 12980 16410
rect 13810 15720 14040 16410
rect 14870 15720 15070 16410
rect 15900 15720 16100 16410
rect 16930 15720 17160 16410
rect 17990 15720 18190 16410
rect 19020 15720 19220 16410
rect 20050 15720 20280 16410
rect 21110 15720 21160 16410
rect 1170 15700 21160 15720
rect 800 15670 21160 15700
rect 9850 14240 10780 14290
rect 9850 13430 9910 14240
rect 10720 13430 10780 14240
rect 9850 9670 10780 13430
rect 10880 14240 11810 14290
rect 10880 13430 10940 14240
rect 11750 13430 11810 14240
rect 10880 9670 11810 13430
rect 11910 14240 12840 14290
rect 11910 13430 11970 14240
rect 12780 13430 12840 14240
rect 11910 9670 12840 13430
rect 12920 14240 13850 14290
rect 12920 13430 12980 14240
rect 13790 13430 13850 14240
rect 12920 9670 13850 13430
rect 13990 11920 14920 15670
rect 15020 11920 15950 15670
rect 16050 11920 16980 15670
rect 17110 11920 18040 15670
rect 18140 11920 19070 15670
rect 19170 11920 20100 15670
rect 20230 11920 21160 15670
rect 13990 11860 21160 11920
rect 13990 11170 14040 11860
rect 14870 11170 15070 11860
rect 15900 11170 16100 11860
rect 16930 11170 17160 11860
rect 17990 11170 18190 11860
rect 19020 11170 19220 11860
rect 20050 11170 20280 11860
rect 21110 11170 21160 11860
rect 13990 11120 21160 11170
rect 200 9640 21160 9670
rect 200 8780 230 9640
rect 570 9610 21160 9640
rect 570 8800 8880 9610
rect 9690 8800 9910 9610
rect 10720 8800 10940 9610
rect 11750 8800 11970 9610
rect 12780 8800 12980 9610
rect 13790 8800 14010 9610
rect 14820 8800 15040 9610
rect 15850 8800 16070 9610
rect 16880 8800 17080 9610
rect 17890 8800 18110 9610
rect 18920 8800 19120 9610
rect 19930 8800 20150 9610
rect 21110 8800 21160 9610
rect 570 8780 21160 8800
rect 200 8750 21160 8780
rect 1400 6890 17060 6920
rect 1400 6030 1430 6890
rect 1770 6870 17060 6890
rect 1770 6060 9930 6870
rect 11200 6060 11430 6870
rect 12240 6060 12460 6870
rect 13270 6060 13660 6870
rect 14930 6060 15160 6870
rect 15970 6060 16190 6870
rect 17000 6060 17060 6870
rect 1770 6030 17060 6060
rect 1400 6000 17060 6030
rect 19180 4170 19330 4200
rect 27200 4170 27600 4190
rect 9840 4140 9940 4160
rect 9840 4070 9850 4140
rect 9930 4070 9940 4140
rect 9840 4050 9940 4070
rect 19180 4070 19200 4170
rect 19310 4070 27220 4170
rect 27580 4070 27600 4170
rect 19180 4040 19330 4070
rect 27200 4050 27600 4070
rect 200 3990 600 4010
rect 200 3880 230 3990
rect 570 3880 600 3990
rect 200 3860 600 3880
rect 800 2860 17060 2890
rect 800 2010 830 2860
rect 1170 2840 17060 2860
rect 1170 2030 9910 2840
rect 11130 2030 11350 2840
rect 12160 2030 12370 2840
rect 13180 2030 13570 2840
rect 14950 2030 15170 2840
rect 15980 2030 16190 2840
rect 17000 2770 17060 2840
rect 27200 2780 27600 2810
rect 17000 2710 24210 2770
rect 17000 2080 23170 2710
rect 23980 2080 24210 2710
rect 27200 2130 27230 2780
rect 27570 2130 27600 2780
rect 27200 2100 27600 2130
rect 17000 2030 24210 2080
rect 1170 2010 17060 2030
rect 800 1980 17060 2010
rect 27200 620 27600 650
rect 27200 340 27230 620
rect 27570 340 27600 620
rect 27200 310 27600 340
<< via3 >>
rect 24520 44430 24600 44560
rect 25620 44430 25700 44560
rect 26170 44430 26250 44560
rect 230 43390 570 44120
rect 12950 43390 13780 44130
rect 13950 43380 14780 44120
rect 15690 43050 15770 43180
rect 830 42290 1170 43030
rect 11740 41800 11820 41880
rect 830 40320 1170 41050
rect 21610 40340 22250 41020
rect 22440 40340 23080 41020
rect 23260 40340 23900 41020
rect 10060 39880 10900 40000
rect 830 38590 1170 39460
rect 10060 38900 10900 39830
rect 27230 38900 27570 39830
rect 10080 37240 10880 38050
rect 12970 36400 13760 37200
rect 13970 36400 14760 37200
rect 17240 35240 17310 35310
rect 22200 35240 22270 35310
rect 1430 32650 1770 33390
rect 830 31770 1170 32510
rect 22440 33250 23080 34060
rect 17240 31230 17310 31300
rect 22260 31230 22330 31300
rect 22440 29170 23080 29980
rect 230 28290 570 29030
rect 1430 26630 1770 27400
rect 27230 23360 27570 24210
rect 830 15700 1170 16440
rect 230 8780 570 9640
rect 1430 6030 1770 6890
rect 9850 4070 9930 4140
rect 27220 4070 27580 4170
rect 230 3880 570 3990
rect 830 2010 1170 2860
rect 27230 2130 27570 2780
rect 27230 340 27570 620
<< mimcap >>
rect 20200 35530 21200 35620
rect 13910 35410 14910 35500
rect 13910 35160 14600 35410
rect 14850 35160 14910 35410
rect 13910 34500 14910 35160
rect 20200 35280 20890 35530
rect 21140 35280 21200 35530
rect 20200 34620 21200 35280
rect 20210 31850 21210 31940
rect 20210 31600 20900 31850
rect 21150 31600 21210 31850
rect 13650 31090 14650 31180
rect 13650 30840 14340 31090
rect 14590 30840 14650 31090
rect 20210 30940 21210 31600
rect 13650 30180 14650 30840
<< mimcapcontact >>
rect 14600 35160 14850 35410
rect 20890 35280 21140 35530
rect 20900 31600 21150 31850
rect 14340 30840 14590 31090
<< metal4 >>
rect 3006 44952 3066 45152
rect 3558 44952 3618 45152
rect 4110 44952 4170 45152
rect 4662 44952 4722 45152
rect 5214 44952 5274 45152
rect 5766 44952 5826 45152
rect 6318 44952 6378 45152
rect 6830 44290 6950 45170
rect 7422 44952 7482 45152
rect 7974 44952 8034 45152
rect 8526 44952 8586 45152
rect 9078 44952 9138 45152
rect 9630 44952 9690 45152
rect 10182 44952 10242 45152
rect 10734 44952 10794 45152
rect 11286 44952 11346 45152
rect 11838 44952 11898 45152
rect 12390 44952 12450 45152
rect 12942 44952 13002 45152
rect 13494 44952 13554 45152
rect 14046 44952 14106 45152
rect 14598 44952 14658 45152
rect 15150 44952 15210 45152
rect 6830 44180 11840 44290
rect 200 44120 600 44160
rect 200 43390 230 44120
rect 570 43390 600 44120
rect 200 29030 600 43390
rect 200 28290 230 29030
rect 570 28290 600 29030
rect 200 9640 600 28290
rect 200 8780 230 9640
rect 570 8780 600 9640
rect 200 3990 600 8780
rect 200 3880 230 3990
rect 570 3880 600 3990
rect 200 1000 600 3880
rect 800 43030 1200 44160
rect 800 42290 830 43030
rect 1170 42290 1200 43030
rect 800 41050 1200 42290
rect 800 40320 830 41050
rect 1170 40320 1200 41050
rect 800 39460 1200 40320
rect 800 38590 830 39460
rect 1170 38590 1200 39460
rect 800 32510 1200 38590
rect 800 31770 830 32510
rect 1170 31770 1200 32510
rect 800 16440 1200 31770
rect 800 15700 830 16440
rect 1170 15700 1200 16440
rect 800 2860 1200 15700
rect 800 2010 830 2860
rect 1170 2010 1200 2860
rect 800 1000 1200 2010
rect 1400 33390 1800 44160
rect 11720 41880 11840 44180
rect 11720 41800 11740 41880
rect 11820 41800 11840 41880
rect 10030 40000 10930 40020
rect 10030 39880 10060 40000
rect 10900 39880 10930 40000
rect 10030 39830 10930 39880
rect 10030 38900 10060 39830
rect 10900 38900 10930 39830
rect 10030 38050 10930 38900
rect 10030 37240 10080 38050
rect 10880 37240 10930 38050
rect 10030 37180 10930 37240
rect 1400 32650 1430 33390
rect 1770 32650 1800 33390
rect 1400 27400 1800 32650
rect 11720 28230 11840 41800
rect 12920 44130 13810 44160
rect 12920 43390 12950 44130
rect 13780 43390 13810 44130
rect 12920 37200 13810 43390
rect 12920 36400 12970 37200
rect 13760 36400 13810 37200
rect 12920 36340 13810 36400
rect 13920 44120 14810 44160
rect 13920 43380 13950 44120
rect 14780 43380 14810 44120
rect 13920 37200 14810 43380
rect 15690 43200 15770 45160
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24520 44580 24600 45160
rect 25086 44952 25146 45152
rect 25620 44580 25710 45160
rect 26170 44580 26260 45160
rect 24500 44560 24620 44580
rect 24500 44430 24520 44560
rect 24600 44430 24620 44560
rect 24500 44410 24620 44430
rect 25600 44560 25720 44580
rect 25600 44430 25620 44560
rect 25700 44430 25720 44560
rect 25600 44410 25720 44430
rect 26150 44560 26270 44580
rect 26150 44430 26170 44560
rect 26250 44430 26270 44560
rect 26150 44410 26270 44430
rect 15670 43180 15790 43200
rect 15670 43050 15690 43180
rect 15770 43050 15790 43180
rect 15670 43030 15790 43050
rect 21560 41020 22300 41080
rect 21560 40340 21610 41020
rect 22250 40340 22300 41020
rect 21560 40290 22300 40340
rect 22390 41020 23130 41080
rect 22390 40340 22440 41020
rect 23080 40340 23130 41020
rect 22390 40290 23130 40340
rect 23210 41020 23950 41080
rect 23210 40340 23260 41020
rect 23900 40340 23950 41020
rect 23210 40290 23950 40340
rect 13920 36400 13970 37200
rect 14760 36400 14810 37200
rect 13920 36340 14810 36400
rect 20860 35530 22290 35560
rect 14570 35410 15350 35440
rect 14570 35160 14600 35410
rect 14850 35330 15350 35410
rect 14850 35310 17330 35330
rect 14850 35240 17240 35310
rect 17310 35240 17330 35310
rect 20860 35280 20890 35530
rect 21140 35310 22290 35530
rect 21140 35280 22200 35310
rect 20860 35260 22200 35280
rect 14850 35220 17330 35240
rect 22180 35240 22200 35260
rect 22270 35240 22290 35310
rect 22180 35220 22290 35240
rect 14850 35160 15350 35220
rect 14570 35140 15350 35160
rect 22440 34120 23080 40290
rect 27200 39830 27600 44160
rect 27200 38900 27230 39830
rect 27570 38900 27600 39830
rect 22390 34060 23130 34120
rect 22390 33250 22440 34060
rect 23080 33250 23130 34060
rect 22390 33190 23130 33250
rect 20870 31850 22350 31880
rect 20870 31600 20900 31850
rect 21150 31600 22350 31850
rect 20870 31580 22350 31600
rect 14710 31300 17330 31320
rect 14710 31230 17240 31300
rect 17310 31230 17330 31300
rect 14710 31210 17330 31230
rect 22240 31300 22350 31580
rect 22240 31230 22260 31300
rect 22330 31230 22350 31300
rect 22240 31210 22350 31230
rect 14710 31120 14880 31210
rect 14310 31090 14880 31120
rect 14310 30840 14340 31090
rect 14590 30840 14880 31090
rect 14310 30820 14880 30840
rect 22440 30040 23080 33190
rect 22390 29980 23130 30040
rect 22390 29170 22440 29980
rect 23080 29170 23130 29980
rect 22390 29110 23130 29170
rect 1400 26630 1430 27400
rect 1770 26630 1800 27400
rect 1400 6890 1800 26630
rect 1400 6030 1430 6890
rect 1770 6030 1800 6890
rect 1400 1000 1800 6030
rect 4930 28130 11840 28230
rect 4930 4160 5070 28130
rect 27200 24210 27600 38900
rect 27200 23360 27230 24210
rect 27570 23360 27600 24210
rect 27200 4170 27600 23360
rect 4930 4140 9940 4160
rect 4930 4070 9850 4140
rect 9930 4070 9940 4140
rect 4930 4050 9940 4070
rect 27200 4070 27220 4170
rect 27580 4070 27600 4170
rect 27200 2780 27600 4070
rect 27200 2130 27230 2780
rect 27570 2130 27600 2780
rect 27200 790 27600 2130
rect 27200 620 27600 650
rect 27200 340 27230 620
rect 27570 340 27600 620
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 200
rect 27200 -10 27600 340
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 1400 1000 1790 44152 1 FreeSans 400 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
