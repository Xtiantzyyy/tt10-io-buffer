VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt10-io-buffer
  CLASS BLOCK ;
  FOREIGN tt10-io-buffer ;
  ORIGIN 0.000 0.000 ;
  SIZE 145.360 BY 225.760 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 6.735000 ;
    PORT
      LAYER met4 ;
        RECT 128.190 224.760 128.490 225.760 ;
    END
  END clk
  PIN ena
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.575000 ;
    PORT
      LAYER met4 ;
        RECT 130.950 224.760 131.250 225.760 ;
    END
  END ena
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 125.430 224.760 125.730 225.760 ;
    END
  END rst_n
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 31.500000 ;
    ANTENNADIFFAREA 157.894989 ;
    PORT
      LAYER met4 ;
        RECT 136.170 0.000 137.070 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 116.850 0.000 117.750 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.530 0.000 98.430 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 78.210 0.000 79.110 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 58.890 0.000 59.790 1.000 ;
    END
  END ua[4]
  PIN ua[5]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.570 0.000 40.470 1.000 ;
    END
  END ua[5]
  PIN ua[6]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.250 0.000 21.150 1.000 ;
    END
  END ua[6]
  PIN ua[7]
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 0.930 0.000 1.830 1.000 ;
    END
  END ua[7]
  PIN ui_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 16.199999 ;
    PORT
      LAYER met4 ;
        RECT 122.670 224.760 122.970 225.760 ;
    END
  END ui_in[0]
  PIN ui_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 119.910 224.760 120.210 225.760 ;
    END
  END ui_in[1]
  PIN ui_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 117.150 224.760 117.450 225.760 ;
    END
  END ui_in[2]
  PIN ui_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 114.390 224.760 114.690 225.760 ;
    END
  END ui_in[3]
  PIN ui_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 111.630 224.760 111.930 225.760 ;
    END
  END ui_in[4]
  PIN ui_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 108.870 224.760 109.170 225.760 ;
    END
  END ui_in[5]
  PIN ui_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 106.110 224.760 106.410 225.760 ;
    END
  END ui_in[6]
  PIN ui_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 103.350 224.760 103.650 225.760 ;
    END
  END ui_in[7]
  PIN uio_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 100.590 224.760 100.890 225.760 ;
    END
  END uio_in[0]
  PIN uio_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 97.830 224.760 98.130 225.760 ;
    END
  END uio_in[1]
  PIN uio_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 95.070 224.760 95.370 225.760 ;
    END
  END uio_in[2]
  PIN uio_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 92.310 224.760 92.610 225.760 ;
    END
  END uio_in[3]
  PIN uio_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 89.550 224.760 89.850 225.760 ;
    END
  END uio_in[4]
  PIN uio_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 86.790 224.760 87.090 225.760 ;
    END
  END uio_in[5]
  PIN uio_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 84.030 224.760 84.330 225.760 ;
    END
  END uio_in[6]
  PIN uio_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 81.270 224.760 81.570 225.760 ;
    END
  END uio_in[7]
  PIN uio_oe[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.150000 ;
    ANTENNADIFFAREA 54.349998 ;
    PORT
      LAYER met4 ;
        RECT 34.350 224.760 34.650 225.760 ;
    END
  END uio_oe[0]
  PIN uio_oe[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 31.590 224.760 31.890 225.760 ;
    END
  END uio_oe[1]
  PIN uio_oe[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 28.830 224.760 29.130 225.760 ;
    END
  END uio_oe[2]
  PIN uio_oe[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 26.070 224.760 26.370 225.760 ;
    END
  END uio_oe[3]
  PIN uio_oe[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 23.310 224.760 23.610 225.760 ;
    END
  END uio_oe[4]
  PIN uio_oe[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 20.550 224.760 20.850 225.760 ;
    END
  END uio_oe[5]
  PIN uio_oe[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 17.790 224.760 18.090 225.760 ;
    END
  END uio_oe[6]
  PIN uio_oe[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 15.030 224.760 15.330 225.760 ;
    END
  END uio_oe[7]
  PIN uio_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 56.430 224.760 56.730 225.760 ;
    END
  END uio_out[0]
  PIN uio_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 53.670 224.760 53.970 225.760 ;
    END
  END uio_out[1]
  PIN uio_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 50.910 224.760 51.210 225.760 ;
    END
  END uio_out[2]
  PIN uio_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 48.150 224.760 48.450 225.760 ;
    END
  END uio_out[3]
  PIN uio_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 45.390 224.760 45.690 225.760 ;
    END
  END uio_out[4]
  PIN uio_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 42.630 224.760 42.930 225.760 ;
    END
  END uio_out[5]
  PIN uio_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 39.870 224.760 40.170 225.760 ;
    END
  END uio_out[6]
  PIN uio_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 37.110 224.760 37.410 225.760 ;
    END
  END uio_out[7]
  PIN uo_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.575000 ;
    PORT
      LAYER met4 ;
        RECT 78.510 224.760 78.810 225.760 ;
    END
  END uo_out[0]
  PIN uo_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 75.750 224.760 76.050 225.760 ;
    END
  END uo_out[1]
  PIN uo_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 72.990 224.760 73.290 225.760 ;
    END
  END uo_out[2]
  PIN uo_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 70.230 224.760 70.530 225.760 ;
    END
  END uo_out[3]
  PIN uo_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 67.470 224.760 67.770 225.760 ;
    END
  END uo_out[4]
  PIN uo_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 64.710 224.760 65.010 225.760 ;
    END
  END uo_out[5]
  PIN uo_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 61.950 224.760 62.250 225.760 ;
    END
  END uo_out[6]
  PIN uo_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 59.190 224.760 59.490 225.760 ;
    END
  END uo_out[7]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  PIN VAPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 7.000 5.000 8.950 220.760 ;
    END
  END VAPWR
  PIN VD
    ANTENNAGATEAREA 31.500000 ;
    ANTENNADIFFAREA 157.894989 ;
    PORT
      LAYER met4 ;
        RECT 136.000 5.000 138.000 220.800 ;
    END
  END VD
  PIN DataP2
    ANTENNAGATEAREA 1.350000 ;
    ANTENNADIFFAREA 1.400000 ;
    PORT
      LAYER li1 ;
        RECT 43.400 176.850 43.800 177.300 ;
    END
  END DataP2
  PIN DataN2
    ANTENNAGATEAREA 3.075000 ;
    ANTENNADIFFAREA 1.400000 ;
    PORT
      LAYER li1 ;
        RECT 56.150 152.750 56.500 153.150 ;
    END
  END DataN2
  OBS
      LAYER nwell ;
        RECT 10.650 21.850 127.250 217.000 ;
      LAYER li1 ;
        RECT 10.650 1.750 129.550 216.800 ;
      LAYER met1 ;
        RECT 1.000 1.650 138.000 220.800 ;
      LAYER met2 ;
        RECT 1.000 1.650 138.000 222.900 ;
      LAYER met3 ;
        RECT 1.000 9.900 138.000 222.900 ;
      LAYER met4 ;
        RECT -6.350 228.650 140.150 228.950 ;
        RECT -6.350 -2.800 -6.050 228.650 ;
        RECT 34.150 225.760 34.750 225.850 ;
        RECT 78.450 225.760 78.850 225.800 ;
        RECT 122.600 225.760 123.000 225.800 ;
        RECT 128.100 225.760 128.550 225.800 ;
        RECT 130.850 225.760 131.300 225.800 ;
        RECT 139.850 225.760 140.150 228.650 ;
        RECT 0.000 224.360 14.630 225.760 ;
        RECT 15.730 224.360 17.390 225.760 ;
        RECT 18.490 224.360 20.150 225.760 ;
        RECT 21.250 224.360 22.910 225.760 ;
        RECT 24.010 224.360 25.670 225.760 ;
        RECT 26.770 224.360 28.430 225.760 ;
        RECT 29.530 224.360 31.190 225.760 ;
        RECT 32.290 224.360 33.950 225.760 ;
        RECT 35.050 224.360 36.710 225.760 ;
        RECT 37.810 224.360 39.470 225.760 ;
        RECT 40.570 224.360 42.230 225.760 ;
        RECT 43.330 224.360 44.990 225.760 ;
        RECT 46.090 224.360 47.750 225.760 ;
        RECT 48.850 224.360 50.510 225.760 ;
        RECT 51.610 224.360 53.270 225.760 ;
        RECT 54.370 224.360 56.030 225.760 ;
        RECT 57.130 224.360 58.790 225.760 ;
        RECT 59.890 224.360 61.550 225.760 ;
        RECT 62.650 224.360 64.310 225.760 ;
        RECT 65.410 224.360 67.070 225.760 ;
        RECT 68.170 224.360 69.830 225.760 ;
        RECT 70.930 224.360 72.590 225.760 ;
        RECT 73.690 224.360 75.350 225.760 ;
        RECT 76.450 224.360 78.110 225.760 ;
        RECT 79.210 224.360 80.870 225.760 ;
        RECT 81.970 224.360 83.630 225.760 ;
        RECT 84.730 224.360 86.390 225.760 ;
        RECT 87.490 224.360 89.150 225.760 ;
        RECT 90.250 224.360 91.910 225.760 ;
        RECT 93.010 224.360 94.670 225.760 ;
        RECT 95.770 224.360 97.430 225.760 ;
        RECT 98.530 224.360 100.190 225.760 ;
        RECT 101.290 224.360 102.950 225.760 ;
        RECT 104.050 224.360 105.710 225.760 ;
        RECT 106.810 224.360 108.470 225.760 ;
        RECT 109.570 224.360 111.230 225.760 ;
        RECT 112.330 224.360 113.990 225.760 ;
        RECT 115.090 224.360 116.750 225.760 ;
        RECT 117.850 224.360 119.510 225.760 ;
        RECT 120.610 224.360 122.270 225.760 ;
        RECT 123.370 224.360 125.030 225.760 ;
        RECT 126.130 224.360 127.790 225.760 ;
        RECT 128.890 224.360 130.550 225.760 ;
        RECT 131.650 224.360 140.150 225.760 ;
        RECT 0.000 221.200 140.150 224.360 ;
        RECT 0.000 221.160 135.600 221.200 ;
        RECT 0.000 4.600 0.600 221.160 ;
        RECT 3.400 4.600 3.600 221.160 ;
        RECT 6.400 4.600 6.600 221.160 ;
        RECT 9.350 4.600 135.600 221.160 ;
        RECT 138.400 4.600 140.150 221.200 ;
        RECT 0.000 1.400 140.150 4.600 ;
        RECT 0.000 0.000 0.530 1.400 ;
        RECT 2.230 0.000 19.850 1.400 ;
        RECT 21.550 0.000 39.170 1.400 ;
        RECT 40.870 0.000 58.490 1.400 ;
        RECT 60.190 0.000 77.810 1.400 ;
        RECT 79.510 0.000 97.130 1.400 ;
        RECT 98.830 0.000 116.450 1.400 ;
        RECT 118.150 0.000 135.770 1.400 ;
        RECT 137.470 0.000 140.150 1.400 ;
        RECT 136.000 -0.050 138.000 0.000 ;
        RECT 139.850 -2.800 140.150 0.000 ;
        RECT -6.350 -3.100 140.150 -2.800 ;
  END
END tt10-io-buffer
END LIBRARY

